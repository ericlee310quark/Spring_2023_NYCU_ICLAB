//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Optimum Application-Specific Integrated System Laboratory
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Spring
//   Lab09  : Online Shopping Platform Simulation
//   Author : Zhi-Ting Dong (yjdzt918.ee11@nycu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.sv
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2023-04)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_OS.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

//================================================================
// parameters & integer
//================================================================
parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
parameter IDNUM   = 256;
integer	Pat_num = 50000;

//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
fvFTdnqk+FHzXcaQqoZOqEYGhUWjxeN8CuvpPBpV8aL1SFmnPx9jUxBKXDO57NBA
4myLioG2O6mbMq6qyBrH+AUETAo8F8G31Qv4WlnqWbhmR3wCOnyQtpkm8+b8G9af
M2DMJHQhl8rlpm7QQ4+WEmk7w9Wab2EZAq13S7OVPsWOigKfzDlh4ClQDfIlSLa+
ro8DrriFmZec9GYf1QeNnvgre+6uLwXeQB/3HiF7iHQbTVLAu8twaiQXmFpo9/fk
Kutfk2s4sPc/OtRKDKYzthJCAHCamXvmVpdo6aqpIP6xp78aFrJNiyCPQu0du37S
UIPGMkDdK1jaSqo3G/eXdw==
//pragma protect end_key_block
//pragma protect digest_block
hn/WZlFyanj8SBkKJPi8tUzlHR8=
//pragma protect end_digest_block
//pragma protect data_block
A6Gbny0Z+fI2qTNwlK20FzXowNd9rT0PWvSzMvcDAjJSrmFOqqgUWJOyQtL4OEC+
ZhH3+iyQKoiIkd2U9ZLt7DDMkBJufdEnWT3YcfItzXe2pkawx2gtQV0rM7nTWM+i
02bYILavK2KhbGrtsVZL0wzSnfWX6wtH/dVJTu1XaC7uZ0ytOoEuOz1DWOuCd9HI
+f7vp2ZTIdEJcOv7GrVBUMUkJ9RzqPh13QXua3o49l+4lVsHgn6PVd3ng6RoVb5W
ZyqmdYVHuupsHv8LyytazTb0WoUz+u/+BrTu6oDeCtyXtF3DJgCr4+1HTfX/5sTm
bEiZeniRwagcLDxv+ETWA5t0vn9sUeWahSL5Q6vGrW+zOkKBHANcgAgzmtiZ3tkv
I5ZU6UJ2Adg6br5zl2AcvYHhB1CBtSGrgjdhYVBzc1/UN7JrGCtxf4QDDyovzupU
1HMJMsH9Dr6rJluA/gKF+APq3dQerke54eeH3Rg53y9PTwIbkID0jk/jPCev/SeO
YL1OpQ9ErdKY3frD71I5ZulXfCTd1XAhVifDtw25P8je6MdzqobCnLani5sYNH72
NgG0fvv/uRCQMAOZB66MSADDlVjyxxAH2/B+03S4JbVkI48aDWXmeVRMZ4ZLYml9
xLUkW8ESRlJSSnQZES2HjWShaXlIEDTTYsF+8mglcwpxg9xIAU8YEY9bMcY5EuxM
0iEfN2dNsNGxTutMF6K4ICu8RZiecajA4rmRB5Pw5YuqFxRV4mZCuCCLQ/bOH92g
pBLwtlJr2dNrRBOp5wQZf+figUVN3AzgDbJdz8wMz5ief4lVTTIG6DmG3lOnBugL
HuF6Gyz9hcXp1llMpl17zDBzPzbxTSDDnrmym0d9rB3BwK58Fz0YP72j42G4hSg2
Yt5Lw+54dg4ujCEq0yUwtZ3VjBIlGDksxI8z2RN0RkYDfmALTTXTDZ2rtNuSwl2j
geZjHTyeLXyTB0HH6TphLZvL8w56Y0bJ+pEfYyGOURNpc/2533/n5z4y5InAJcXu
Hsai6i7OA6DwIBjFHS88Ows5yPz7i+VlpIIRjUaiNateh6lDB3khhzAvUeq2cQ07
Sn/uRC0YYHlMhqyInjmwLwj/JqurIUvpmMRK/VmB/k4jc6wW6U/NYw1f/xGqmF47
3uWyl3SUCrrWYEcB7NmmqgbQL7WTeUEC0h+5J4ouSPVvvLQTTnD/h2A3YVpbNRlr
IK7tKbf+cBi5btjkWrrmvchgU8YLcn3q9zKr1HhyWdASxUuSpdBG9YPBzQUFoH/o
2V/xDL9RT3R1nNSjJRML/5ImwIUGk8gX+6zyUNNzn6pbV0mAejdWP6k8pBssa3zQ
A14K/GEA2Hmti8nJ1KYVQKJ4ujjZtO23JefOjVq/gVhh/PmX3hgoQvWdqeL0tMNV
NNoy54yR51FwTwubL/3n0po0OPiF+JPkaSZS0OolLBvtZwIYClD7uL0Tme0a9XeA
Q1P3/DD87mCHAWLpfnCQxLrfTnqjVaPnHLqthPpoFZS7A+QMKj7besZe8M+aptvQ
k5Ya+nXaQ/RHyBKhxkUAiy+0p4RzxmEnJ0e9+8jYYablUAOw0NF9EPNLjFeJ5Ece
yDt+biaWpLOymHlbp8M6jF0Vgs92WSkk9nlkRNVyOQH5e1+1FnmfMTiojhTgiWhA
h6czfqZA7jc0BG4GH77/Iz8QE7ta3Z4DMr98IS/7rHEe95e5tZqi3aXRQbCoOWtu
utcV3j9SgWBw9mI78+F/0nFOIEjLFV/pFlwBmRKScII9wLD6k+hORzG62K8YwWGL
sYEA5xZ3Mv0SgFhQWDZu5jB6ebFBSrk+E67ojH1r7tRSNAs0pWT4wCKy0BNyWs/i
wud81HfKoB1IVYHKx/WCRqMTTSUWwjh8IEjML/+k787LINzXaX+tSzTLbMorXVro
qB1xw2eQjg32G16qugryZ9CpAz5yP2FL4wUya7dqayI3IUsYPI6SMs+WxGcm19Ol
7XkW8PEBknmB5H1pcRRSsYDpYOu1Y/4v2vgMWVIAV4DmcmSKgDxfJyrPlFn1EOHz
q/+fGNnXBsh71ii6E4cBvR9Z34Pw9MMLhZBjq3IOoGjKD0H+chSWryLe7sQvTWVa
U6nT43VVHLGAOYPBMWUNX50haT8efspWRWUapwHmiWJC9/gMRnSH5wd9Zzr8w1Rv
IW0JgTHhOmJmaVX9WBoimkCtZFj/d8Ln6EsALkD0F+lLepEvuV/bjK7bdBizlC57
jtpHRq1ZIkVZhBAHsBprSosGmFEiAR5CffM/NYd3PGH/j+g2c/tic24Pdxn+MxPa
PJJvGH//KfEiV9T4pgH9XS6/7+vsAvrPhXquCEcwP8eHfb1ZAi657dBCeDmZACWy
tL6P196s0hHMzLiOIF2otqtK7/IS/U49L8UNN+ACFffgCLegM35uxzZeie4lscrW
Zys6QvZHmBGov5Vf/ikuoc3slgGcwmYsLdzCBSVDij2TuC9u7TXKIWy6yRVUUEoF
1apGCbf2T6AKAUKUEeWgYFV8Plfj9V5Lvh+Fc5KEGTyod+NFBt0+DfYvExPoXBrv
A2SqLWPKGr9YD0MMS4cQysRPCCB1aLI34cLrUjlSs6JbiJLvc1df1MgmFCpaEG3P
99CvSJxZSPGj9wV3K3kiNrtxHkRq1CnBQp6/DKm+Q/9klMEhbsjxZVnXl1bDjocP
8kit6M9q+UY9RmJCbeWXYO+tmJ471tACRWtH6NLQ2TRMTXObbGmDCnCb6WANSc7E
TFR3ozjiSfXyJzYmfugUDIQEXpOuDQqtrlMye+kDu9gPOiioIv0YlD6QcdPqj1Wf
SoDPOsJnBpwtGOFGLBf2MahtUdXp73kKvc1WgiLi73pv4eNXqJTxhykM2mwUC+MZ
nKdimlmfZoAas9PSekfQWusEqN8LRHvYLIEVl1zC7OBb8lpP0aHTYKbDk9nrb4lK
oPMZztwGUD4SEq1A9aHV9wgwD3Ua6A/el8waWOaEg/YpE5Pkie+fu2zK/smCWuiR
pM4sTLU7gZPlanTNU8lWyvhsLVSh1DLrE5biS7VawHKY1hFovhE3HOkscm+pomZy
QCsX9YQMZphCLDohmHaX6Dwg1TBMQA3KgMUO3UGE4FFQCGaBbmKrcZRrPUD69zyB
a/5v4650SY+j4qqBfQBHy8yxCNAms5WaikLCujePBPZRfI8ARa3sH9vLIE4+/VK+
gOmj9LMV76dNjuKKP5z6T2owPf3RsdXh9qdEo492nlkJR0idMlx/L1/jJhjKt9Cs
L+8KBORCdP/gxFwPTqYCeA+PW7A15eRD6TLnG1EmuBvcUL0m6ABEzLzkBlc/9We6
N+Ze8KvS3loZ3RwdHA9vfuBIjI1eyOJ+N28iFCRbW46jdATQmytySjOCmX+/4ShZ
kH+upNzJNGPSgtvb9z8lmv1bLNY8I3NSe8XqN58jRxY5etLPUECwolJ0olUgZH3n
cr4AiJwNgJoCL4TqFdInquNg9WENFjJ3fXNvpPRgwKTXQKvXSeIMjzqCFxdJKxK/
orxAdzbdYt33KEVsZr/zSzDbj0jANn8VPSiARu4q9k8rGSuMrDekZYTKP1RgHXp+
r3lIpw0McPy2gHcky7giAtq+RBro7SLpOV/mB6hWJh1/thTibvgmjIaKwZ1cD6hR
WnKn5DQrxnDbkrGYXVChNaXN6dPo3LVJ6+VPXh5vX956EphkB1eYbSJBKeTmDTMg
PvgfXKEHlB9gNNqRziVt++zETefFL09tUWDIijWpr1zk/x4x04YlQ2RqMcQW0bEw
ZitVMHkkwZKgFQCuGBjowJSThcLdP+EjaVAj2wzDWU2MuIlnOhqYdJgTI9gfCSvE
akXRrmht0Rwq5AsuUrhmQnsv5iZ7VQRBD3hpayGe8wg8kP2IuEO5eW6rIKcSyTIG
4XA4NcNSL62g1q0mugaN2qYJ6Qs0ZSGN97+/VkGDhu1tXQtaSYS0nsI3SbqeQplT
bf+oph9csFjE6BPt1sz0BfrrzqCrm5EL785UqSE6dkzAknuPcf4AQQS9+lrr56Ib
kpxg2kUWviZE0ZxO+y5+XnkHU8tCZJ2oA+GuCG8wdrR7cA/7ZcwNl5u3gdcfGR3l
pn0NPFTlk6PijBxxN90lrcG+gEeysCwVc32wtcAowPqF3aRkc7sI55UuON9+Pm5N
I8gvlJiMuMzZuMESf1niks1sM3ldJjakkAklWvsNoXxNatpf0flCZKZKgdTT6pXH
PJ6h1BrgB0e9HebqrZqqKG1oKSONblEKXKcBp8CBRXbFuypQOxfj15skFqfvXFNp
+nd8+YLOmp2bvPrtyPgb7iGxrImima1a6j3H8Oc2cAL0zekVBdOsfjgnX1wIbVhg
z1BvYYS/BllAQsBPumK2t/xUDkcWOcPIHrvikyAxX0W/qRP0mgjT3R6mZrLXZbof
r3PIj3RGcO+M258QphhVWNHSKyZHt9bJyulvlw3UasyVHlluVNr4SHRB+CVRn4YO
fEWQL/YVNaH2UWsgEWFEblj0OUe4w8sL4DQbQDNm7xAoOdlpXshfoGWNdBJTC7Im
P2UobDeBbMm2slNN9+04L6/2nfIW+k4P1dbdxCxdxyIUn3e9BIbrAIGuQV0T4J/c
FuavMh89APNn6nfKhIhKYqAUodnbujWe2Y+8TKO3ee0n8xqTj4EohKlrUb1ucy/H
Zkdg+VItLhGRhMx741L04plXh6FRTSLuRHD1cFGXYBKm41nmvIVPL8xEhXa04Ryb
2ZCvmdJmUFMTKl0MQj3v3JjDdSKtK2sNCA0QLcXZ0klt8aX7p4Cu4sboZKne57pJ
EzbBGc0tp58LwFxRbi9IuHTAyY9cZ7wydA18eBINxJcL+3mc4pYKxeCtORqPyBFR
rL+g5FiaOhCn4WBIoLdI5ApVSbZbz+GKuyslY1AFiBl/sKZFC4Ma4WFCL3hlU0vr
ORZ7hHit5iDp4ylOylJFrOz3tLrWS4zp+r2//l5KqAFA50TYuiYC338T3nzoAap7
vdUzZAVywtCtF0qtjPBcf++TQcj+Xzn0u4n2c9KwDintvFmEPd+qmG+blXKYgnPT
vNzKLXD3JUvZXFItP/mUoR3wzN0GtJ2XIIMqNb4xVbIh1a22/YU6zCBnsxMYuXqs
QW9rv05l/THvBCmHTHeoqQdahOa46UyTD3RL8QWZiQztHYyEQx5atgMtTCK1cdsz
a23vhF96kNBQjFxKdkXAkEwqMdxQzSuzM+iE0TBdzlXS9N2/V5bilvYrySvT8kVf
D2fRZKr6W7RneS+a7zCCd6hOCDn7ENLuoY2AwWPBX05Nc/V1iE3CtYD4Pt9PnKmL
wggszwROsfGWMZyAwTwNJOUtOsQgNa4zvAuRcQcDerJrZtiUBLHy7/LOOl5lhgLk
E49I2wk92CwEZCcIADjo32Iz5kcP98xebxTlZ8zGBIYlB5WsA3Qk9QGpyrs+iyGn
bJMDsAMs+7O6fGOiChbqQD1ixE5btQO+GSalA0UG0+/mcvuklIkDzv3Pblg2uJ+y
Ns3LoAi61tK+JGY1DxelRh4Bq3FJW2Nu8kPXV6oT1xlxsk0NotZ8J6BQ7n/spA27
awGcau2EBEmuuWRd38LyAaFzLDhGY7SAX9eE63+QzOPCd50OYGRIMrJBsIinEp1h
M9+vvB4+/JJ5y/rRFxPIsDVA6SQcbDgCGsOndQaZrLozFfd1qKXtFcyMaYmlvPmF
ie2GTtIwDgAU1VXwZKHuzb3gILpM33d3+uIBBKlNi6uGoTtmsHWkmBGNEDbaMKeJ
R04NiY5/O8DDWokMCMmkmr5LssNVk+Td/l/AeUNd8bHlr1ZBI3I6YtSRIJNcea+t
DePWsfiAf8Xg2B64W2yVdaQrknUXg1WgQ/w4oFzWltL2cPDQg4/AnKlF3dyMkX7j
k1bFOsqwMq0obBcf2c3r9aRZditrR6F4DCLzwmonr86e9zEplr4ANrUuzkP5u0gt
XHmUtmfKrzixp33Eg7lPyQ9Q1EPR49/iHM3uuu6AbW++yyGppNITqX9qoVUpv1+h
BrpSAOu65fZxVl8vDI5vymkRY52PgXdZgakIQGSYwo1Bd1X6/xfKSh45BfHmDpm0
Kdmv2eWja/7aSAzDVgICM2yvwqWaTKJZ/7S6LShhqsS++nbP1/yTipT96LsWVJZZ
TIy5jEud/utUV2BQf4+Xmdcc6Kh3lin9z/YO1z4f9LWUdZnWLpisSuIS6C29Q+4p
fatNW30qooNo1Ru5LTOETWMJcJapcoTqOM5rRpOR/oreSI6GT+ElKLub3A3yMv9S
glsoA2Im7qwHOPKbraPOpH+P1bGp6C5tCFx8GcXDdk5hYTgFJL4slTbraX2rtUsG
OLbZQzt2rS7P7K52Tk4MQBIRf1fxIZKlSFTDEueptS6KzYoQt0wX8Il2Nsj0hdp0
j23h3gbVYj439nUVp9BL6APXlY7/nI8lxSP42rbDN9uxHXcehWuNmOTLCX1gHAbW
g7kgJJjhsm4ppD2ezgTzlOuZ8EQJb2pNTjU2LjlIVlyeC+YfKX06NHBlIk6a6fzV
uarQouGfZy1lz432mzdm4kHU45S8fGJ5wy1OcXQnBb3/HZ4ESDX2d/WayaFskQ0V
YYrczYfgQi2weAQ7hcvOXNAy6c7O7DOrLBN6nzXvQ7vFuhFBNK6wRWfnqy+qZxjD
3TzuCNuNAemme1yZrvHbYJNbUA+Iedm3LaR9m6uNvcOkBL+CXXqUOyZBOGThFC2z
DGtVebTNs13EDJTQzkHm0bUWWwqSLBZckvFDqRbjyBipmzh0s0LaUlk95MacWrqJ
tsqWbmLJX7b8cRoGDn0GMBmaHYXmKKma8Ph1PcbfNwuuQBTpG058aMXQKJjXedPH
itP0FIRmNHJp4ez3yTgdLF5p39O46X9dhvkwU6Sc4aW6tQFB50Fh2GB+3P3x7VLL
cFp2LCnQF9tFRwIsfYOc9siVP5YOlj55/jVX6Q6ypk6JdLkDANZZgGyOlRUjyDvi
3vrJ5ebm3noeywfifeM0nXo5A1M+l3RO9NPpLdjX4SQnBNg06v5e8ylH53Fv3yuP
HydQrOj/5U0KJ3tXAxqIHi9QSn+hJClu5dMWXMped6FSpB/a5VfQdVTdnJzBe5Cy
TNL0gO0F0PQb4wndLZgJz5L0DAmhRYK+hO7Zs6wPW7HKaqc3qnMbAvGdEFzbs+AX
5KCTBpr5NKE+IkN1uuMwVEV1yQ4Z+MN3N5rS1JY4sODvxWTNmDGVmtlrCawv/1po
e2PxsTI3Xr1sfKixzynvNYkFALR3TVbEm9YsLMh0LG6mPQt4yx2npHg/Is+qX87o
IUzZpFzn3shlw2QYbrzHgANCPWW4n9I5NlPdb+Aoo2CaUprytPGxTMJlyyzC3d3s
15t1bqCVqzYjgNvidzqr4qQKMnQ5EAPec5CjUACNCITyJUACaOMUQWAnWTWerHFN
CszxL3SrvaHCqii/c/hAxIaAvtA2coDYLA0t1U0QXnftY2wpIx9mJjBeDF386oMr
teG50uLUUcYCx7VWpr7COZ1fb+/6Cte/T2ALZ+w04TJ6XLd+SlO6zESxYl/MSlrW
+JxXVWpWa8vAT9hvt5Q8MT8bHiHflaIMXrK0IV6esknJDhzEv7H4rCsF6mHh4VQw
ld+Haa6rd/dbMSnZj2/MQXz9PMeX5bbFp7m2LEkJHCrOUBTUiGnJuiFlxK9OzAD/
C1Vhg0chnrglIc9yx42rdTQy2B51z23tNEB1T15UO4I96NRKXld5zWexFykp+lXc
wzcVp0eDpRf+p8n97I4dS8HjgqZ8HYWKZvfHzIn1QZaY+b4MTs6ur+rHLCzqm+VV
JZ4pXgGDq7uWcN8BYih3B817CYE306QTOB6Ox0depDO4DK78dh1q2vl0mmDJ9cw4
wLkhLX91usd3bawGXvop1jNNJzgcbISm6PVA+CXrm5cQrO0dzXRwYTcy2RZOk5Kf
LnsKTa9hrgeREZg+i9hTTFoHdI0OyLHLoln1WgfZCDKi6RqrmvbGQHM7mDnuYD45
UaK6z24CoAK7tt2mNl1gVCgs2yxHl7fWzD537Ym/lzpltNkb7GVgAdSwd38lAjfq
lHkpIeKj9QYGYx1Cl+H/YMtObwQQ/yhDTF0dPlB0SZ5BarkZ8virI8RVjnu2F7aI
bC2PM/GzSLl+HID1WoSVJNhKah2DP89Rp38/trenzV611vZY/7PrPyWqonAKl15R
+4lujvr6P7jc7NyUi+ZQ+vjtx73npTqXQxVGY4pYyIhNi0KrHjARix1oEsK9ABpc
/spHP4OH6jLx7JV0AlRWJTYHdYJYjuuAmgMrFJa8rNoSeTkqXQjsz1hA5kAQ8gvn
dWBiIiWpLuoskhkZZtzwBg0NtqZAmlpojCgfL8lgZmdNnn93EY7Kd8izxO8ufHXU
DMSYy0wcuA1VMWYjRDRRfdwBqFWP5YU/6Ww0VLy9XaXmFUobMTxKjo3HnHwljMr3
ZZTchSKBkyjloEUEudIXRAnqmUFHccBLIiXoXg7CnGzQVnZ0SlwOGHnodyTG3WSW
AkbS49OjjoKtBqPmdZFdLXBVzyAsshqlTwpVyGIp1+3ghbx5Rh3n8xXSAxE0y9I2
w3tDLwgPwMqadRMOp9X+3M/bwEEWWIfpsAdLQ1dz7SJsgr0rNmTTf06DKF/ZOXFr
pmamddQ9/0QZG7HPxBQgmY7WTpmUT8pEiXR3nqFlsOxFig6YhnY1cJWnSXFlESe4
tJh9LNRo4yOeC9J46NvgZXHT64cH1vO8aVlNOkQhTBabzHEfTt7HGZDa8hzoMUQg
VwXqzbI1VbglMPdSArbqoDmaFgMAM4xVs/3fQWzafr/nZ6kjbcPPbQz9fQZhaLH6
tAmSDR3d+mc/3mQanFNlQiE2I+yw2sOZR+uWSAAhfADQlkPaLUj2M4zIUYmrzHSu
i0PrtJIkcKbMgBj4ESI4ToqrMXs10c02mSxTqcPoxFl9rhMOYf1FIPqO8mjf38eM
P4uUNki9T1UepBPB2jckkYE5vETNeHpAE656lIf3ARWSEbX2skNSTdrvYp8lJSqb
hCeIhDy0diIynsAjjmcq2mV2DWKCROx5VDoD4KlN3rQzXhds+UqMbF7X24z+qjL6
+d7reLtuzXr7dXiY7MGTkplRtu9M+aPowmh4bkJ9ZQvq+e8vrH4NULNVYFDVdJxQ
TSo+59/X/35vbp0r+rA6j5x7FmpiYLV2omYbVH0FjX4SWsCDu1rGGrAmQ/O1tm0k
GW+D6+xnX7zTk3E3Aq+tm1R0m1YUWEq2Vp0T7+SZDnPwe7J2kTNpsWsWAez+6fUb
6Un6rLHg4T15jCK53Bz+UdV4dd77SHkcShecc8XyGEF3m5mM9IfWF196+IKN7ZDy
QKtAL+k2QbcKB/qJsUTXySgWtPl2wEZ062xiOKSl0g9HMbIggA6TbGjdRJRpmxSY
Gt3B6cgrmFFFC+MxHPQf1JryolPHVhoO9lnWg02FSw0uT82EMEEkoppuIWuHJDKA
SL/tIoRREVuVfhj9eAMB+nDnfrCJ/iz4d+yOiLcacsk/sY+Rg2BB4khwGqeSlylX
bH+ExOq9c5CXC+tk3ANsxCc2d85nJy38R1NOFdpiF1tyJZv7EUOtFb9U2jq28lNh
gQvgnfHfJeQtlSgsrZVCdA08OczQxKqkRJRIDez9ZQv7baiDvIGOVXJB1N5aoGBd
Yw2v8bffRmJeMx2Z6Iuk9R9bPyDhvCYDarnPMHdQYJrgsmnNkjCpsJDgWFC6xN6j
w5CCxWVOwIWK++IjBoIZbIgMEPx6xw8jm9bLJMkT32lBEMU+hrnOSRyDtZ/jrd3d
Kjy/Sh+nGXVHWZj6OxZphdpfCCmVnkOkw6tniEh0ZQxHPQftMi5NhvsdVv8qYAS+
0KATJ5htzQMq2OlxeNtRGxL5niHPE1LowxsUSySxNKQZLqH7O0brsRDm3UBlbb/Y
vRDLncnK07YDPSf+INGYLxejSyEcX3TsCk08FuvACflztod8KaA2XVF2NOnTH3M6
Dt7mgQEQVeSAyL9Q4idJFS7Dph7o9cRHQfCzcXI70/eiWp4p/Stk0pHyiro0kgXE
KAJlyIdoj2tyKzkd8unHJEATGlQjdrdAvl8ralM0j2on3/ct0bWxmFatSwMHGz0z
m1IDmvcjMecdIkaLxw+kwpvjZNzaGTQ36IVgceMvK2ogrXxC8c+RDimx3o/EmD6s
Tx72YyhA5oa50e5llqO6D1CTIVBsgS5xW+XGESsAEd7Dx6dO1uyP5ObgG8H5pNrG
d8LjcBIsnL/JUjI/TqkA3K8vxex89YaF5KhH7y9PFC78mhd4tOozsjVBqQyofBa8
Jnmd4xZ9G8LQCvh4VKFZ/yeKPYRdn/DyXJbUm3yEMLNsk/D/esoxFFbwbqEjqI8I
SuEQDSSU9Yf1a8uVWSUcm6udZ7uzgG1LgI1qd1XNBZc3zPVbWO8HPudsIsub5P1C
p7UVrfiwjPDkRjS1BAf95kfCOWxBRmcNsz0+PsnuvG3/GuF4VHGLJdPiSSbee0na
zy8XMSOL4Cfc7Pt49mz6e0WO2w51Hnx8MwoFMgotGRFTUvfzVm1jICUIkCYdb5TU
uvyuKaCpqTuNkruRjb5Tx7VrNC3/hznZqx7k9LHvc29i58+V0TujFoRjc430ptMF
i5BHrXkp3qjRxB7MOTaMEfg1baOlYAhYQ4U2+RFgXGEpBb/Z5/6EZ+n6/nmZUMRd
H0mF7KKEow9fpk3LFlnYgy8YL9mJIOjvn+c/EgqeIlcd5qmC44Tcrp3HKXYUCsds
nPm308HFP5rKH46OjdVI/HOuhRGEF++6QA9NFXLShN0UuKBCoSKaDywPIJmpXMRF
7VZs41ChOAJhp71HO+7oix7rrjiz+W9SSboj2mUHZZ/yfVoXyCfKsOKEkKiPr1uG
JO++n+IXGk7V8o891n4vLhHckCHsJMqywk9Q1RqNgggyM48aCWhr1iswd/ZXo/Ev
Z3fYmIpNavgbUBUzFOPaa/JQr7vO+8Znir0KY5BqW7Da2R+nvAR+FbZAgQtHhlfD
ORaae9fvOALiGgYIefn67ipgaWZ6nRwiCmlp1aqpv37cMwPKYhAk5qTGyI/mwYx0
y/2FREBVDPYHA96EdYZXAUrJTHF/8g/Yaq5j3EzYC82gSfAhPqQn5VitfFQ7e9or
pqgnWc74hGXMZTGXh5IJYpYZ9kaxoIbtgEpjcCGHNb1JOKJtL0xcJ+6BzQLelVOS
d1VXlD+9A3m/YBhsuAzwZPqb5+oM7zmByqFmcYfxaPHFgBswuDo1ErRF1Xg7kVAZ
r/A2wTecUsxjyBGo5ODURlNbmXiYR7tw0mGQ4PFWJXqZCybLI5DTuI0jy7Sq9dzp
URnTYWZ7asLAuLAVH1ZL7WoqkWSugitPOKp1AbEHopvSFpbMd5LiyJcKRt3JIE4w
VPKu7RFTrgDwzACbuSsC5RV4qXDvxkrSocoQT+Uw3kLfMaLYFEvcUpEUr9kW8xmP
+4qhPqQHOcoS0UvobU92ceD57XmENdFlVpd9dEKGigId7BjEz8aaa1XqXNrz7A85
aDX6eZAoPAaJd6SGOq7ylBcJJY5pNziVqXSLlueAg0wnm+B20xHuGyf2oHqExgmx
Rm6AFNPUC87I7BmLEWCxWCF3oL5p8L49ZsIQxntT4GqkgpoDVX/NMXHMPWsNucdY
M0BvHiiTyg/VWEYdGv1T/WsIELOxI6FMCoo1bKef0vPjGF2M4omu/7NIkzVLAARS
vYRCdsTag+xV98qC2pFSdu/m/PA+vZwnq2hstfrfhYKQuqrSSHEQRLQnIP2PDPSu
x3ZVweA0RGytmxB5zs96QGgsB9cz+5tNZ/ve7Uxm2x55likvtgTcBYyB15fGZffC
fFpziKYT/4njczrreHeh0xn3NRGjQDbBBKEe6IzQl18cCXTXuIa/qJJKq3b0+0Sq
hjPdXF0HeCWHQP4xwV9f+xGeULBTAeOhfKPDRB+RSOIkFS6N46tY/u7OGygD36BZ
j00xbE2ToA7Q7SyWIdtr/ARupGtY+wFhLvV8Axt30xaFpONWsuif1ILuJWMe1s8X
Bp+1iiYlV6DWTOpZ2bDs5QEW12mfb2DI6XOPqm7IfviWRmMYzLKMUmMsSjdpuOnO
7L87JzCMuQtG+DB/fIReRskBtP7XsXxXS9TDkw8nqxzwaVkx4BTe5PXGzKGUhxvK
mZyHkUBMvSqb1+lKmP1v7SAWgtW7d2qs2jBVScfwWV2/edaqUetJ4jBHbHPT/Lke
ywptOQOWUVtJfCeR9YK5P2Za+VoCeMxLCcEwpeBelbtDXcBZani+MSyeblqB9vfd
k20g1GLEIHwZC82ZBey74L+GWRDpQlZwSILvrUQVv0yH4iDyWqu4uYxApTx9Ih/H
ktJIZWGSWrCx0VQR9PV0dm87IYMoswhxr0EQ4BMoZ1D7XDe5DVJpwXJ4aehZtMUZ
VRFsnDY9bdkJYMg1jVhC3IrDyii6CfOmNLgrKM+CBgtrrBNFvGN03OgQEqcUIrgW
WpnT9/Og/2LxkD2ItEKnr5e/9sgKDLxQpzeo5GWnDDF+1b6hyljA2vftkrCJ2Q7O
7svPwBTSHF78j7O03JyXbyhymHHp+Y++a2rpKl5UY2pdIAOSrqG+s2SHGXQI++li
N4QG3DO/tNURCuFjFQo64RZtIlS05l9YqYBOff6u14UoW6UWqT37kkMaCtBGxBak
sIrgFVvKTEFNnnr4X6S/cX7h4hqAdob9PZDUgnNGkqQf/0gdjtnITpsBC7dIRdpk
mPypkjvk6LYOa2kJo2s4pb71KhyRv4BKkDq079/3coeHV3eRQ1s5qYxAiUm/+i/3
SESIY1woaDGORE9/K1/9UEUwyMfuNubYBnAuFwVQrFBckWSVemq4N0y426M0w1AZ
X5x4PqwYRMNXRJlA88+1hUFmMA6u/x61rD/I2W6noTeKcFV8unQ2bu/DWcolxDCQ
bdrw7ftGpT46xRG3mIwpGdLIecKbIXf6jrIGjhzSWrgiZjBCJsmk74GjlmDWR/EW
zx21vytCJY4AIXH5BAImvpdpNtBPQkGZn1qXTIGn+pmLx9TL9gaYtlR6vGcBQLau
TUidTxRx/zsN6Nb3dHmFTKb3hSQDs/k3D1xXEH8o4iIaVG/5KrEq1CUQ1qLK+gDV
vnQynEQGMwrXE4b3GgkJCRQMI6f/nD1qQjPsV/PtTku2Wdzdkmaf7fMOZMbNbxfO
+KPycaeKIxyyzoxJcfhqEkrIcKzrVxBO4zLyIJDMQCWNkdXJUhp803Arz2xgSyB1
U8Za/ghQhrADdNgY09aVH/iTyV3N1YNUEB3yXR6BEKkK4/xf3LNHq8F9fSKsKf4o
FnPO5ynLMJdSU6eHAO3QmR3bbGkYfe1p9aUzTNJdCtEVRLwDspynf/Vqzxcl7Xkv
kH+45ml3BPjj7dqG5LtryEZSzdnN1yg5ypTPuYwvPVXVIOl5HahRBrcL9ZKbYMaY
pEbF+Lfm0vIZdqWVnTtwR3TQ3Si6ReZHhr9M7QtKdO064mLQvs8rj2cWii5jUfSp
daRm8cHldRq/5B/NN3SHJbhuS9xC3McDOqSifDw+TTpS6h+qejyNqxD8+1XgqAw0
6TtRUcDskCVos0iajdlCg/dZnbfBAbB43V5geqCrGyWmsEwS8k1Dcv4xgmxkx5TX
CArmDeIg4UfXAK0sg3+tCIlrt8klSvblkSF+/iYMT60Un8vRdZQ/p8WGzRj40ef5
9WN6MOTmVyinNHwtAjJYPjXaFXr0zFQiVNZM2www/N991SOczaVywKRGlA/QSAsQ
x2f70p+JViEDyh28EOphUvCvtboJOrWZAtYoXlxtRy4kMVM6C/zu0HDTnjz6xCPd
4GgCcF7gKjW25moUSOeT0GmIlhsxMprAkwrDvtmZbbY4jSOEhc/rlTq6yr5kTS/3
I/mDChQbJ+gIqujKmh4Axydeaw2+aAyaAmzNSYdh49nnpuEzDhqn8JpKD/2bqB/M
cFeMIm/S0Elzml4ZjsnrIJly3jXOtJOOX6GNO/UPr05guGSaZyM9aKNUGebsNchT
JXcE99g/whznbFj7ocwXBO/vHZrJm64aMTTiE7IvDv5BMUFOQDlRFeOBx+C0UHm7
5b9ki7s/2uP3FeW4PN1DbQidbU9l1/tKHU/UdAn7tE/h6pX6k/7b/wRcCjk61F+f
8QIB5QH7l1eprzZTvv7VmciEhw4BheugGaj50i54t1YlWPCggQozm22ky1aMoAU1
Uc2jXXWkqKUQcIDp3KcVnjLPi7It+j4X0oz4Pr6I6oxUMCjKl7xQC8h0vBcXXy5T
vjEG5Rmd2fwCHOfx9/KlBxQuEDbDKlk8MhXVgJQAkHEcbuhlU9vbd+HBAL2963h6
KZ3SaslrEFD3A2kShsvmwnZjnd5wjsPn0SPvUO5TlUjDF6GsGCW+cDw3vlMJTgBu
cd0Kyhb4YCzd/B2bwEyGu8B8Ho+8nRJwXx0agYGS5NHv+pKkPsw8bDts/TdI9q14
D5wVwV8nGCCBkwHqDfwv1zyd5oz6u5KM5VKyn8pv+8xvwdw79RdxrI39KDEhNBxc
DMzFM+u/3BERTa+wDRPWe+fTx3I0nv7Htgb7nC6CKxsS263FL+ocwtITWfqhx7EI
VXDMJlWKaLRRswTeUz67VdQBx1xki/qIXRMWVrYA+wMO+eD9peMuMFCG+h8OJ3on
T1tsfoVyPXU3rJlJxPBbh50wZJBtyVJn5TgHssH4GisM2sG7IP13cY7zjQUi4TeA
VYUV17glrmQLPq2axd5M7GhL3N7qfCPacNkJstibxIw2165DSw77MpKTyRblZkQE
zsM0Hr3Qoce47YdEWndCyCr1oBWIwW6vujobaHaCpEfroIqmgjSEcXLVqrdSMG0B
9JAhSv5TleI466kqeVneHfcuh3D/Xqf10VBhlEQgg7LznlaCti8r0Mn1fxb0YvHW
fpaBkp2ghKUuJ7rLIs142m9Y1NzDwQ6NSk/Ai1cR9AbhIcJmgs8O1jlf2x2RuyyL
3IbogVYQ2vizV30Uj244AweFfeOnhtmdv8Kb71TdFEb4/vIedsmL0pTMD664RfZv
lZa77eJXKvemp4LxLnmDW+S86OKdUaT5w9I6sWm64j5Lwl96QJqtv78jShikZboc
cJF6uB1efCmaypT+4e12FUpcRaLJy8QvlxZQRahsyHJwgV09c4it2KfyFyUS8mp4
X11+0QN+kwLl7DMnpyIfsoN6OHzyGHY/aTfStBLLOhUOBtdorg5hOMPAooAFGncU
RRGu/y1iKF4bnhTpAUo9oswQJ5Oyc/S0p74JBKhADArQmSb0LXOgQH/kenbVgIZU
E0G4wv2QOV5ZtzAJa5H+AuF6GNOeuKTo9yCGk7Dogp301X7qMt4sJSiPfmbbpJwT
4WxlPIz4NDRMusivo0T2LSmGxs8dLs1AcNNwjyUcqyzA4R0LsUCe6a6bD5PZx97a
Tm5JQ17XOHvqftDgXodg/CP1EVldEsUFP9eLw1SAUCdwBWTEuO/KuSwPVQatpCvb
B1gzi//CSABhTiDNzt5aJLSp8l4t2PC7DOqQx28gXXeZT8OMckggWUdlBuc8Cb/9
bdhjvslW3ecleXHPfhMzLCukrIx3HzGgV0WQ+5wbpMQDgul5ScImm0Aq4p8vC6OZ
Szx9ERaMsb8IxTgsl7VPScxzZQyGazg4GqrjiPU3PknHYl05SbtrF7nUVMaTdQ97
RaAFS7BL89n0MODY/MjjRVG/33dZ/fVbtTiaX7AttDpu1eVNZk2Vw1XCp//m03Rc
SyNT38Om4OX8nFzm1kv7W8pfoAHhIhaMKjA47oAgLZYn6mVC1S5FR9XJVjLYY6jm
UGIAuTDVS9mpEHE4L/AbjFN49r5DV492LujWnPz50j4H718KDSelAR3r/Vkka52x
Qfr/InQ/iJadMAwmguMXAdLiMBGJZPcVDu1fnzrmG/t1ZuDy55jxyICcqKqgdPcy
X8/qcd6QWFsnn9S5OwyGBwLMl5UAoIKoNYSILpxPIpgN+cgpl37ydsR+W2xiqRgC
phAbYBOV4+sZCMdDu5Xlmo/0qOVWOFQjjTETH2ByhFkjy4eVUaVesth6thT5c4Xg
cvs6mjgvWFckylY6bLobvAQzvDIGaMtsgyARuMUelRAlMRsqs47WStJG16Z1Mubc
o+sosKL2+vAIqn1PQTXuLoxIz1eWAlHBdqcCkdLPRY2Q5aP8RHUaFJjwCl0gAD+9
L38/BZ+dsWi1246fHvNZTHfBzjX2px4YjPYKmT8hf/mfyGw6/BFJqVqZp8PPgfcA
2l0Cto3zXD24NDLvKAYaYwbOAzDaiWtU8pkcVouFvIjp8Io93pWQnnh95HUchv8F
6BMo82EHETu+rwom+v48Lx4CdvtGf5FJvB2SBmdnM9fuGUU0Iklfgb2Oz7Imo8AS
l3metYs1w5WOnOGZzM5Lf1iQLL0PBJ5dcp42AlVpP8PVNe4553rLIrrMSp5CLjDj
2oMuusiw6v0TlWcI0dZA6RWvX079bLCNPFL6VmC7secs7WBj4bxpRuefUAtv/sBB
jo4+lVQM4cNKChfoWIz8h0G8v8MSQVmjeVfuEdGpiWdIRWHeJXmhR3EElfCONXxQ
Ddl5J5kJH27V+Pedcr8Eq4P3CfuOBxZJQ6Z03+Z/VX7raumvu5/w2Bxk2Tsn6xHY
bWsgXLBdT9vSPNEyJbWfxXz6B1c8WZNAvnDrNUifBTUbdZnCRKeoPy6eycv1Uczr
txDzMWoBfDhum0RZAMrmbWsR/LqnynLxFiX/4g7otVZyeO9WLnmQ7yl/dVhBSica
8G50MSrUcTb9heBxTjDbKcIQ3Sfr+qTz//iVseFH1YxRNFE9b7Q/qeFE3KHqQ2nL
MlgrjVb5UA0cn+5FtVK3cUUBjazwA2z+C3hUr6N6WIn8VNyHA97piI/br1xIA7mR
B+EaT1pk5XurGoRg3b9tENOuZ8OxIBwBAe8Vsh2eoGTHY3nqWeZEM9n9b2Xh0IAg
n+NIN/U2FIE9KZhzW3Se4+2bfjOSRe5echyEumHYsBet18mvoMV68cdl8jgOJLIH
ZotXpuFaQTf9W2TTm3C3FZmRBHhdJN3X1pYp+aqJeHq98pVtffvu+sqd+2pnsrbB
877umrasVc0u2PNNkYvoQUC8CA+oII7NjewL5/ca5KActjiwwj8KacBoulRXdkgc
SaTT8zmYAuJZQ6luDi4C+cJecbakvCub9FacicpRAFU+3lTRR39bEphsg4dv1hyO
uH+SYBLv8j9h0QUhFoTmiySDqE0n1zbsEPymoCnis19Gemy3Wuq1Z1VexvMqJ0qZ
aTWaNHsXFNkColbZ4kXFV7g+3hmi2Xp0T+6VLqU/cfJK+oyi75czVCAouvlqQhxk
RoMWD2qk5V+q/cGpkMsm6mP5JwnP/u0UnOWrgyrkM+k5lZDNt+rmzibafuNUcC0H
+u9U38Sgs85i+kTQAwGxD2k0zcQvjp+VNt2+cpABVy7L+QcjPmO8kk9/UIxUzRNB
8j04CYnq9sHXjzI0ul4LH2cmmcRqXWibI+BWkJe5Reazw4LW/fxF8eOj28oMwUk/
9qy8tQsQ4+/pzRUT+kMMMd0kFfPYeMRK24+E1yfqZYCV0PnztYAVkGZol8XORCYz
NYx+MlPRVwOEd8YtQKfouF22FWfcm4YfOoKbCvdsMZ/C6ynQua3mW6PAP9gvsR7N
c+L345bXVOSdL0i7fk4CUZedvDZP7o8wMtHtAdKfTUf8Mhi50lZONQ6zzCVmHW5c
cqB1ImN6XXQOM26TlZh+0PR6IjFuFsdcDU9hQ9GVZiv7ys+I61XC5aUhaTlnrUMv
37h508+2zUiv2A6NNIO1jg8Vu48UHPTgkfM6pB1sMqbsZNmphfv1B7DAdE7inVV7
zi+DaeuccbOZue2zzy6s8rrO/dol9ifKSwi8Xz4Mk0v3hm23ABkWPyvV4oqLQN3p
FxtFragB8ihXnq+c54CdWHk31/0of+FGXVq93tUjfqOFlFkyma2Ylxzmt45OhdkM
8b35fmJLIymacTuRu3d5IjbTvF4IYSM0Ks1+nvkNld+zNW46ZpEWS5VlUS0/R4op
oD6hbzjcBPn3pAz3x4Lp06XkwuB46jO4bBP4TAtfk1U9ocxHeQZRmIZvQZY52N4+
C120bwAZaMr2SCSMI2UQmg/VVffZQZ9jbuS7mqWw5EzSeVTCesicXAWsSJpjRdaN
WsAJUGMhQvFxxXVLp8ifFTWXkyDaWA9hegpbW49qHzAGXpWEVAIxuz7y4BdhlhWe
gnzNJ2xbgWjUSGEuGH06sjuhDvpzsgsdn/VAsdyjAqbUCUHvJecCwIIMtVd7Kpgu
+HMzLiojM/WezgzgFsQJukqhsc3Vhwkz1sVqxZVZhE2ZmiIkDmUcYVqw/g587hpo
HUmkUL9ahn9WwKf++s8hY4OGCf5BZnbvO1tRDlx/a9S1t/xPkc5DEdn9TcxgAgnw
3UP9LycSbaKgeLqsgAsz3fBjBsH1xrhzNFFq9BqnQMyuw37HAV6k2X3wc8naBF4j
K+LBKtNhJrhgvKSJx0oq+d/8jTiaQsy39KiHKZGYjIHzU2+NXHvTrnz+WlDA5O8a
DwlETLr+0CRZ4n0mxGuC8XQ5E9UA2sDxyD+7a3DBsppFjcOgQlO++0Q+KzG7YTh0
O6KQZw7Z8ADFG7QJZ6TbCweVhtROmhYzEyChUVmcEm9tf9Z1Kxo7mUFKE4sHK1Qb
tdChG8UvNESgu3w/v+7gV//gNrITtKP1QZWvYB+rnOPzSU/02c12ANK8A4MJUzT1
on/+CKwcZe06CpsiwNKtYgiAKeHl/2RcYd3lk8GVr4xaQo3GmQ1TgPxkmcNh94r3
gzAiIvCdL0yr/rUMxVC6X2ObKvamkl84Am8ro+YQDxjFQmF3E1BDypxeXyD39w+X
czxk4mTeLH5+VbuZS2dKWsSQZ8mijL+SQqpcNhN1KDF1rDW1iKxlwppbSfIeR04p
7+SenkyiizGabMWjzrxyA1SbWCFe6wwhK8OCa6vj68goT1dMwH8meZmeiZhZK0kS
twwmiNM6INJlYFPk7jjtw+//WIPOqEMkS+H+6c7SqEAtlhTi5r+TMSRIiMklwR5v
DMe7v43zke1v3LVtbtfQ4Kyeg8uU+7XRRFXEzdWl7msiOIe7i6ZxEvtLgowOcUCs
KTfNi/acWKCCibtT4rotey3VNMXHOQ8b3w8OfgJdxT+/f0KEbenG3reaRa34GrAC
R29ab7UnH4R+zChaMLBxRZVj1pJKMZfXG8xGbzYJy5fkzc2HZXc2PK6fmncmv92m
hzPr+IOHCioyciXwyUdX92D3vmJU4bm/BaIoxOB/ISsgjpsSzK8G8EuhEW6VSNc4
aW4jkIDGCOi0H7bIyy6fWhvyYTe+CWIapX1Ga4DVyS21dr1ljpnTYwL+ogWUfZEk
X27His9um4+Y6Wwl0y23vb8bvMPL/81WOM6vTTT2poIXqf/qNT+i82sdAnfBudm6
9L+YysPCM0z6AmXJ1wlhhz27Zo/ctctjUMOifGdqcFJSuEj61iyMqMfNvjqx8ESC
xUIY2Vtdn9VQdAGz2KxCxgGMihvpwh61SWFjfSyD35RWhNa4UzY3aPvqpMoGU065
jRzH4HMTLiRSjDx4BT+UIQJDN4ImVRflkoidvNhlsBM6TEGfeMfBkvijEpXLCHGV
K+fYMLtLRyw5wn+iVOF1K5pRUHxTCR70UTO36J9ntWOvK0c7cf8wnSXcosCl1mJO
cj7HKOYkc/lcNJJsM9dw0QaDEb5En587Nhg/6+ZvNZfrEAvo40VtwhJK/azg9/GC
YxJxNMMrLuElMpo7fZZ5YRp0+ORHSqVD8OtCqk5THHorbJKJejn8412g86lo+WgO
6Vcp/oCiCwj8sNKUdvta7hixjGVNADepm0nZ0TVujvGge1e9Oen4AvxTpEA/s8yJ
0kdHNm5SXegNXjuoiDJ0lCtK734dcW9aSZVRx9Y78TFh9rgDtOoAzSYV0TmmCWC5
gZlzeNPzIWzncSfUrCMGXNep+3HDpIlzgynp1tEx+07qun0P17Sb0kEF+aStM0cQ
7A+gLrXWcII8sSOxflhjrlYuT+eFLBgtaco6NLbMfXLu9YqVvGQvOzUgxexeV4oy
Zmx8Jsh0I9YfzbsjikItiRutxA4c+frhQLQ3A/PEp2ZHOVi/2zUUG1ee/YKVcy58
7u6utGYu+k1qn0LaSKqn4WEipUw3KJsMP8jjvHxVgmiFlX0xb0SA8z3krGBLUJi6
XwAou7fBjJ14ycQIfXJmkKPMVFV3Df1//0hoZDI6cGeZjo6TW5qkc2QSB96t3/69
XjvczI9LfyV3XkFy7HGjZMOMY8YLT5zCugWPvk7es/NEXUE6r8ge9fYeb/gZZZxu
K0t+fCTaShCDizqPbzurTEex/Yo/ia5mHlXiqTSYJl+J16SycAkzaWyI0jWerDDK
/bl5sv6GzluSLH0/u2A+kjqeNQKtYjxSz9ixEODMW3Q5iOax/zLnBEbzmifGAWI8
TF6hYy30BnywteRTCEjIZalhFg5PkSC+kIU7Kco325RcLwPVx4VzCrnSNzlHUtOT
Da1miU2wdeU1bmAKCL5Tt/gw9yr+WWYoSHpuPYQ7sn4FAixz5LqrAk8zppU561T1
Rv2zL3QAQL/rBqy/RIksdYW47MRoOLmKeRhiMAzWkHUJfgT/aC8SzLc4ntcdszAd
kY875u88OHn0u76UEISR+0O1ZZGairJPL64ZrJYlucipaNIV5t6MZ/mUYzq7iD7T
3Ex51nU23ef7qX6R+CATqL3vXig6aLqm0XaF+DQGF2cQE3KD39In6SOjK/R4ZIw9
vtWjh3n1oIaWDlVkvy0KMBIwq5hcLS4J4pibWA0yH7ZQDQuZU7KlLF3qS1W1uetg
530C0TSNkdU/6pCVFEoxLEHwT51R/tIo5knUMGFXq4OdVlHDqWJ3Wljz7zjeJ93t
5SKSsXfrio7faierlVqQvGRqLM+YaGFNdymr5MQziDKakjsM6khOCA7R45enu+5L
l5qGUrV/zTTlv4OeS3k2JapnWLMJP0dR1TskCxL2B58BibJZtJnDpWKPJh+LZkTo
t6C5AWSPdm1iX7winK3nvg4nzQuE9PQPlIUYYQLezZjt8c5MBM2quBR9FmX+NN6A
WLjTiPMAxMQMIMlbCwDEnnasyuu6X7GXArRCwQxJB/ILqeZbMb63oiYcO+mxH4H/
kMFzkM4m7mWN79uUfyXuWNF0etkBLcToky50hUVqjhQTyUXEaEJYLquM9vKBJjyH
CZRkepPcyBD8CCtAoQ7KVLej85VMH9DtJ7Hoh47KJ7JeGD/hJd6MRQ3ei7I4e5z6
VNAezVIzGqqsyJSZvb49iv9U0EqLv4z52X/PrTigf/cJf/HyWKozNJCw8ke+P42i
4YRzg9DxrOTmmb1iwHMb0kU1y7dX3tJ5+gPEluMcelqoTqcd+tWsa9WTX4ZEeinm
H0onR0HOXf10dbRmXz25htHO5O76GFDW+fuorahfZfKYoDOvmsBRVqdHkaDJYGk3
BIoVgqoX4o1I7MVxU6ilJDUVnkd8XP41K4HDIqgMiYWpS6eYEZEgqmTiDIiB98uu
ZOe4Saf++VOK0/nQpMg1duIk/0g8bi1yebYRsl2NHcafc73zlwJqrDqOy+41gaKS
x4RWUdS9qqJmdExpbvUGhg7t2NTd9dg0BA5YhCZJkdcZyb8vX2nDowIPAP5A1TRy
rjvCYgyLf52AYsgslJIMkEJCwGmqjElNu5XzAS+TSzFZaBuCIpSgLmRGlz+whhwT
3i+kz0XDas6g5bTakwwo6Kmaomg7K6LYXN9FTyLqqCCdfFK0WG9JnPILh1vhF8EZ
8nn0zY0kZvzBzxKkyMTnF8kmdSRYngkgmZeuVMlxNJtK6LAZwptEUwHPfwmMjmA2
Kgbky2gx3wTBohl4Ed2urtqkFk7Oy+3AHpcayfQ5exzsp+aej+2jE1HN+Ep8mRZX
bSzPSkrwl2hE9kEimxuXkXjr9KS0sLJ4NtDAJK+O2TUUfGY5ssgGYsdSaWlUI46x
s4AJe3kWCoMkE8iZpL0M+3uaBOtvyjUY49RqYvPrHPd5RbnbMX9C3RWjg0RNP94X
/KGnvuJjAraOOZe90VpzlDZC2nLdq4CwGpqbRhgNJNm2LbTeQ+KP/2bAzcmalDY4
WbTxq16VVMFpJCFmau/HUyuYVWu9tJKjl9QEo8zU1+ZFhwVaaB47cnOpuVe6Y11Z
zCiMv0oMQed8HM34UY2WIWplJ7avAcZQ6x1hizQrSPes9HvFy1fe4zYE3hIU8QpM
xWIXkWZlaF2EMq7PLPPRq9DtCVUkFfbpS3ybEui2sxfAUCnSWaomMkJ0HTwkg5tQ
cUnixcP/A2cp/2/exhzJ/XxNT4BQWdFERnWypA+mEjJfmlPeqmtP3QlIE/FpHk+Z
M7NwFKbR3/ZJ2PNCIRpW/i2Fo2ifjp1YwB7yMiUpf9dKJJ8iF/eMQaHU/xavIY/L
nAByzewCr74PEHRF7solK2gV+lmySXg1L+WCYh7g0qPY05TQAMRDOjZE6EP2ghpP
kXUChsx5Q8RRxjnDC2+JBnPXjeF3IjndXdLnkmBk4ELUxCDXfk46QWP9yiMbiJMm
h2amgFZFQF6DwZhkFYs8I50JHHQERwUAGszhqjp9LZNZbCXtfISJpqBC6hIQ1Kkh
qb21ET96/aZQhG0hFDCBu06JsnSxt1z0ei9yzzw406lvN/1KuslYQrD9E79Y0A97
fH2wATpJElsfG8UCVb9l3wWU2u020NTXQsK5/LD6gn64D/g89ldk3tCDY5jdct9z
kHksX64cQVjeUMhMC50lWQ0iZ+RnU56zDFC9HJ4IKAFv1fvFwIMO+ik8O1/7XiUi
t84LaMc8ZYkX957vXfECN5BrDbmlCEk8/fvNOov3CTNUY5rgbNyFRhmd9kaj/8zN
dgHrn+WqKCwBOO8m4I95OEL0sb5HRuTlYZjYYM0pQXQu6NtA3Yw9TC3Mwl83ThoT
t/6ZEwAqjbtGYu8nebAWpAP78hOGNOGtT8+zSuvSU8b80MEW/GIzZtrkux4OEW9L
l8tCta+CfApSobE3q7HiWRPhBz1SxMftV4uuvFD6Q9cNiBcEL+5iixlg/5bfGCNm
DeRcqnOpKMramaCavDvoqnE57hQSEgudjyiM8QKIAnoL134zETIFTfl7uN58IXVY
5O+BV14gvdi+e44dLC2ygU1jrVNyODkEk87qjjppsyMpmHim+Fiq+64mFgy0sgNQ
JD0BjM+uOqy3GNr5i01CKMNjK7Cc5n48Mu8wjw0qeiFQ9K79EnNWezzytU7ZdhGB
llrOOMiBeGvSO8gZ0QJIoPIQkUKvBmH+fzVoZFlB8Sqdy5ghYm6LjA6yHuSNMW8y
ijNi+g8ja6BtiYtFRUmiSkAvSAJsTzNWKkouzciWF+AxQsl84n54ZxsBFRPn6q4O
6kSR3Fyak4vBIZiSfgNM2yAGFhCquBe9FIKhHGQPuvcwKFxBxD8uh2Kr2qx0TpBU
dUiNDvQYCxEt6j/tTaNbKXaVNll5t1biPDzimxa1qD8g0XaCWu3sm8HYvpK+TZnf
AzTrqLtnLBcq5t2fBPoXCjgukFUZanVesTmEZGGFLcR93xS8m0nzx4mR0QsAFQpV
ohFdso8Pf0bPgkYdmUvIZF8VQ6a/tq/z5J37DECp8QNz3e1LfhMBMr+JckP+Vx0x
xaRviHC0Sb173EGNbFpYZZYIw2QSectXgt1eg4wlR3If5gQukyUl+zZ7V0iwvKtc
dy7EJ8kMtQOQQTcdEe+dP/tkh7dC55RaPPW7W7fPnG434t0ZKNw2ZddJsB43eqyP
mJKuT8C8oDfn2pPU8XliG2Lz2vHv8bnKd3hszzvlbPgmRUePsDw0e1auPW60OiwV
MlxqQPsw/oJXr9bUy2HoRLTnxa/jwJQIqVcYVK9FKj8apcJeKmPQYN3k9WwbCO+C
UNxHO+GRTxMgN4ZRNeK383/QhK/R6c2cBc2BV3WPpfIDACd9wSHsg47Oj5Beui6n
rFZrFbAMepsfE0Ku4vL9scpmW0nxQx+oE8bKXsfYpd+8jAq/OBOdmfukIceqicfu
dn7rqfIkVtKoIVHTfo+mmRK3FfCQd2QNsAyo8ZFRQIospY8icoslSD6zueFBg/Es
z3rFwwZODH309N9ZE+diKOoIzRBvJD52gv/1m/8M1C2mChL/AhgmFW72wNv47OFp
SsBjmaET8yNpNiPME399vUgtzrGgCLd+37i4GNd1QIQK/rBdyWqhTWEb5hoEI23H
CiC7ZcC95OVdLZKlligjlOBngl4mC//VQnywupvivLWLSyakm01syJw2fzE77bMF
J0lZ2vFduRXuT/WdWmB7BYCkO5Rjg/x7F8U9kAAQanBSmPuTv6SlbTmtcLodOuxj
9kF3amiiohRu0Op9Vnqn0IOY6ecFYFovO7kbbYzvBLaNAP1670uqb9nmVjJxmpHR
2a3Po0PFI2BuVm+HTZ1gUnRVIhFjLTa3bqKBJe4SpUEAPuVJN+dUC9pLuxsQZdfq
xCpcLXhOdFZt0k9Hs/OEun8emcn/zxJkYe6YXgqxzZHE6Cpc0DTuEVj2k8f0Sr9O
VcQPtqAkdxYFcmbFfPN1pf5dNRw16gawN6n/Vj3KUUXEEGs3NZlqyUK+Y6j5kfCH
DZLJ1WUvMtVynY0UXCM73f7T52pop8EeziSIRFdhs+aMNfnkxBRR1lHCyEQUSkuD
OyI48oZPQBMQRF9+u5Glyh+o/7Rzan3sqhtPPGqnTKvBPzkQv7d9awJeNyeON1Xm
gb+wkHX+fpcBpqzeSHsxOtow/LnPSz5QRoWvqVLYep8IbEHx4Rwa/am3aqoYZJQM
c6FhlA9Ti7tov+dqld50O8mbsdxkChXKz4DayWermUrYqLnuBOh896FoL7Fsob+h
c8FcC/LBzQtIOcI7Jh9VlJXQ4kSt2rJXn+zqHyqg0dPHHwoS7tif1ZSNKwC5QuuV
5K1VF/BttxxyyHZmJYF37uhsZERnQB5WfdmkWMmKfdd0bWVovwryFlw9DGD6YeMm
2OfKk7WAJJQyhNAHJ3NZFsJfhEKfMmnkb8RmLi/nvbH9rwlUACLgElKka035ImjU
3B/5effltoD1e4H9N5A4B+j6k4+b5GyDKCRH72T4+a+d8dKPlPgsmeDlB/r8DkSm
XQULxwG16ehgnRZ6NQKGfSjmr9KdjNr5Ydu1G3k8rOtfEQ8XkyCV/B+tzIk65QHt
H3B6zWQIHajVoJJsONvQqvZ8nwQx2gYAA8XKCwc6dObk3QdOCFIYImysTIblRkja
yjdT95KBu1/kbECKAf/rZx8TrXp71QQ39vJmZhew4souznrw8kY0kH6cGGk9wurs
cqX7XGCpUOLTRMsd3egZFWCmDx5qwkBOwD9hxbw12bPqx6lLZn9UOLyKqxKy8I8p
HKQsxqsbLOxhXJJdyAjHxYzLNCVkJJ1ytnEzzD0T2/dHEd/jX2jf0cWmhc6hXIkX
6FSFPKMRykP8T48ct08zt+xuDW+qS4J0bAZ7emTgVCc61h9IUJ1u6Zl7DanrGJ/O
RRDMh11shpDwHH9yMeffxMpKXAHMnPbYnskbblp6gJhTkK20NVLC7yXP4YKptZUR
ndAgyk7ECgpYyLHe26KeAkpb87vdTjgKw5Hz2SeFIuMsFt7FULhUmOwDpOfiEhR/
OQDN70eTWi/z3JKGI/xeXZwrHHLCspnxo5YZnEKPJfDo8tQTMxRLMpfoBSH10Ywu
1ih5xyqq6wrcOXVmWPySwLaMp5sgneiZFVMh7DMDsY6Cedpgq+cvLn06l0BeNqh+
NncFfxpU+28xPcoomSgRg+TXIpooYYK6HIsuAfJagJSAt1fRZkkUpyOXdxP5R5XO
KUk8oz2/CbeV7saIvi+ZPEWeIjN0KNugVI2Qj/a5eriUJBK5rwuW/tkeMmPyA6Sx
NzTR3BG+Ju0uN3lvlTMd39/D7rtuteR/8PjoUfrdW8fNzdhaA/YJEoRgwyTQm9Qq
yGeKMkEwA/f13pN34Z7wM6qwAKoROgEicSq2fs7uTQr1oLgZJwLI1watJ61afu14
O6LcLb0kkpjrB4WvVATRZwZQXUreRQiDr8T3JxXDnqkTU6VH6DivXnRpwZ8ZcFuw
zRwjbestEL0gHZKtS5PAp+DP5HFp3gn3nrMP92GQ2R8Hll3VyN78BJV7P0RCJERB
X0TRhq9pbsYRr3JJMw+jXv1bclV99YRbH4Z83KSBE189fI9FQaO/sQjz/UCcYc7E
gz4ywJ5O0OmmxarsbfpV1PtHSCcgBtWwl8gvuJo5FAg5MJZUf4gOALK/l9goKMBo
0GdsBJkqCc7xdPzITtQunQQ4/lp7fuKxLWb0TPa+rmppOgwm8/epA8DgvX1Zzqj3
8aTR6Br67JekSjpo26GzUj1Qgx0c02kwKeDusJmKehDA3QXo9V252xIs2Knzc1On
a0J+nrn+ZTS0HkYeF3qxqOwvEsreSkGlEQV51ReBhDhDANhhdmzBD6CbmkXvkTEx
qKxyB0Sta7SvQFjswHq+L3FnZHGIwc0bhkB13TCpHxsy7dsQy+0Q8Vhy+zWKZlPM
FbiNqtuejbre7fvCxJQXS4wF6HEae1GyFN9Y9XFlFz5W53mEvBF8Ljmka26pTF9J
+eTP0UvXgVm7Sa7iagnvi5/T8YVtEgn5CU3k5O7AOIaLh6qVELBKxuNW3TPAOtZi
jr0kvG3MNtvCzkpCSekcbwCBBMVd0kf9rdF+ARFM1emr4J9tlzT35fr4yYFw6Bfe
T+/qvFPyEY3kKuvxcU4Z+MXbhAIGWPvjqqOYqpmIp7aBDyJt2p4e3PTBdG/VbX/g
ELGGNwQNMpFVbTb8vUUshsDZlXlhRkvEa0idrBNzwSqi2KzFK8lwPqMHBBWM0B17
Hng2KIAR2oAK1hvweLYAMCKEWEwwlkPrj+y9vTj3oSSK7SneYhRdtuB8IqDW+VKM
vGa0VgtmkmhvC8XB2AqpJNrea/GrITfYxX2gt+AueGVFJ/PVtdCwijvEMuqEsF1L
fVZFpzD8Hux2SlEnviFGDkvz9yhGJ5hSGzOcPReJVZgLuUcL2OwzXgl7ULl3J5qk
itF6J2wPqHpboSakoZ6vXWxGaHtWLCCLJzMSNz3SQU8CQ0D78io+hU4uOjPUsAms
l9lhPU0ezJ/jd5Et5k2BCxPjOLHT3kG3F8lIMog18KhH6HVojB5fNBa6NMQk53EM
8WUbUI1fBPVJ4KHJF33RfmWQ9VM+J8YsfA6oUQgWD71yf4fdg5pjM4trp35PvkPi
vzQFBUEikR1s1axZJrAB5Zwsww6iVFYVvDQodVLTlHUnFULCkA/spV9kwFnN3JPO
wpDLrWbo9Ial0EXdqd6DWKxs/I5eaFohiFwS7YmqSImfpn5UG+3bed4OAVndXRJ8
6ck8EIVIHARDSeLojvu9clcj5sSHe9BcLsMHnYHOPSvKP3FfWXQ73Se+VcdQFZ1I
hEvcIzeDHeNQQ3W+ndnjv4/+40RUblP301RJVD/csT+ggAELE8olv3xF4MpN9581
dzPYPjS4ePBke0yD5DzH647IpQ8HAU1z9AbK7mkVa2nrvzRB0Bo9zB/BvqECiUcN
LC1HtuMypvkDSesOrq/xBY6azI3rXjAt/Ou5nNlEt7opitmLbjvgNbAeS3yPVe45
VgP9faqtmo2+V3oewGU1nwK6H5tl/m2M56FsnrUqCjMy8nEm6gf9wGaiMxUvkbo3
9j5Pyt8MyoKTitGZQSqfJ6u4MGMILR6dxJHVp0W7RneoAL8r5TozvmihmH1XI1wp
tA0N0qPN0xu1jOUtGKa0XdF7B4+i0BfCGn4MBv57KHWlcBdys47v6ST9zOukPMxp
QX2qUAgsYJVfCm7uEH0Qxxiq+lvoLu4s2/4jRso/CxpXHtbr68wAT039X+A49J9T
4pZkxPHtwSznEl+PYbSCC2+8JIroaSJ1G7uPVaSp5qJBhn/d0Izdk6gOMYUL/2pr
EsDNoPzAX8wtyZFavwK7RdFg2aUtIVcPVX6oUbj3LhhTxMdDIDnqYz0NzoZ20TcJ
F/S55g9+0NMOZ9efCD76H9FeDr3VGQRaD5vzHm8xu/7Ysq7kKxwOjgwZuPldAo8l
NxeAGGHl9BMubDoeggl2PxnzO3OvBZUpJiUnbHYYTp7b/NS8W5CtF24ZuCnyGNS4
CNZgpRP0QpEER0WGiecHxYK7ytSpGdzl6XlcHJokz0vJBVhKT5UPdPnoqn/aTu/J
pmOH127qzIixdnEWkEv/NdZD/qVXkykTgUesEs0F8buHjt19UsLVO6raEYOZsn3Y
7db9A/j1yPS7/3TbLQysM3XsvNS18z6V5Vk4h+BQ1AUEW+Uge8SjMblzA5GtiyV7
B2owCLlFsWcegMcuqazhMuDvPgoUQNbbNjXezX+nFXnTPDS67k1+v6v8A3VCE27U
5ZxYSOoBEZmiS6Ad9MniB6aSOSER+pd2ohe2TRG1M97QmwpaxQ9D5gyP5vxkp1AG
ViiDcOZAkzIip4fpPVGjFHNyVMJOu+hRtGeGYjMnLaCpImt/rqXkB+yQkoHwNkvq
xgESl0ZnCRExUUqI5GTHjb+yTJK5UUqRq1LNQKgQnqDCOuZewHAfRT1tR7PZzb+v
6VIMUP/EAGKePegd9sOpTbmFrsv4rO/Qg1yRsQ3T9ob6qdTHcnpjcr8y2dY1ZtE8
SlppOOhP5gL26wkTbm2rgiwNIHSU3ohVPmCuaXbywKsyscbdH9piQIVtyPU5dyPr
nkYkk5ph0JCzxulqh2ve5gNmPj/iXJECfoFX6cdQbsHI2mAsjuLTKcHA+0fnFwTE
zFtrH1bDMe9HkzXMl0ubaPKOqWByupYyvInQ+H5EDL+5KlAYzoxIXbzxLoBUtFvo
7OKVL0RAlWVxWkVAfsRrO2HwWnfpzyFpBBgllrUdBtrwqLMI+VLTAdLI6ynl6LJt
knhzfUL4fRVtOuRRE7zvIzbh0d6nRBei3hN6IR+zdyYmlIB9J6lrah6xwuufQN0r
6rAH2QUv/CEdhXGL4d9T5uqBtWDPx29dxlaMYopf82QdzIc/fSxZQkoCz5HIVtm3
nTCA8aLS9Lv8OraC5htC6vWr4i4IM9H3cUFI0FuG8IZzPJFEz8czQXVw3B8HiBIs
orAeNGg15ygYnoZpr85UEWdKPzd4t43hBiER24HG2njXjTGHIn8a0EhZ4MCr7op7
PjaeS6hOU3HJ2LHH8riDLhGbYhG8Vpfzk/xRzQ9bysehyVOqsOp1jZT8I+/e1Y81
qhc0LpuldsEnQADFHaK4kaZsWeGxBme3AVINNNgowGNcucMRPF9w/jLzR6wQs4fN
HzNaS8AfBZBlPRvrV5vu2GG7bJi3Z/kQ6PA60Wi5bOwUen8jUXFhiDIAVBYw5nOt
e5g8lyPncn20rgIpEU+p6J9ZECBWqFNHRUPPg+NK4ZoJu11b2my1cZ0mDla8ZAFM
amUZ/5PAantGwLexmO8+nDH1YFlyzfm73rFmJZX+mOn2VlD2rZVwHJNAJZUTgULD
7slGFSd9fCaqn/cTpnMnrN/ZiziNAG03bPNjlTmFzc0UNdwVw2oHQ7NZAS8eJEk8
3JlM9MCBcpPy3IREWkqwavsyMbcjvx3DVg7oQH+SlHqOpeusFB3nPWWlL+inCHKg
AXC78rG7rTYa/ZEcgGF8YSYGc4jsILu0zIv4/qxr+FB9UaAhjXyE8IMgive4GXGN
7nrAPT+iZFduEM6qPAKo5XhRJ5JI5+qLxOStfiTmIQCbiZcotV/Js2y+kUx774nx
HqJ43qCo54H8tOlaJ1hfbIVRHlacLXsq91e+2gV/0Mzg67uogPJRWGK3it3f4OD7
1uDg4DiZZUjBKiSuWp68VL7aE26L7upIRT+kjP0VU3nCMgpw8Bws4ZB2t2qO9qGp
TJn4ZmKB6ZRZzPjIhzmnzhQiacA3EwfVbPHICMSgUinit+90Zr9lq7D9tEhYt1jU
44d+5aijlau6C6d0puS8ZNK2ryenSw9bI+UQVnvwDqVuYdR31J68EmkZJhGrMWav
SoLx4wfXlWElrFyOCz4rprPjCl8M8qnoB/o8LyEw9PSOA1OMv6JdxWAiYS/P+k61
gIvCWRTkJxAfA/J1F3x/kGN/SYYPixob7hQ3j3tHvAvJF7jZYSruSMyGmP/HLpxU
Vfd84g2gP/BEmBpW2g1XBw0pmlhO0zbuuTZOKCwnyKkm/QroQjOhdwo0nZJk7Vz8
yRoWAkZkchRieY9QPdeH2JFgxOz6WqwF3Map/UQGBOS9Eznx4lQV8uSehykrDO3y
hTNMUI8kj+5Pj5tphINr4Va7rRSfOYa9AkW6zFqH7Z53PGWZllY1PB++12yOEwmR
Yo7+FgZmeuocmpw+lTTQgXvVBio5hdhu5iUfAGWUIW9zEVgTiTW0eYMnzCAOeKtm
VrsGKeo5S2oclwFbIDt2ajIga3aXiVchKAMTGe9TsdL8vJ5CMCYyRDjs0tZAF5vn
eEm/eDoPjeBRrabFFrOraoiKJAMXG5dzkzO0puAjIhPwxS4Ev16I17+7mGLxzkI8
tLWRMhClEat4A5GEiWt1NXTNU8x8xhL1gygji95YTpcZ/Ha5UoWyDDsbJWVGVKyW
pe6P97wwPf/AORij4V6JU3PAxdfzUluSYcPevXqYXQ4PgoZR1DveUcPLpdtp+qEz
/BHJgEbcOQql6G6BXFcd4k/MEPt1eAjfW5H0Qr2D/e8ojep2JjxaRGnycLQyrHJl
GsoV2M22WLuPRndb+mfQeAyh3yKvqcD32ki63pF2KBSHsYoG8urbdAvLiB7cugMO
09rZnCizDL9aZsRM+r19Da/fkFF0CE5lLidU44F6J/lTblUOP1yjP41THQrbMHTj
W6tj43nXmzEJUm8ahH4G8J8ZIaIWxYGmDFvn1vI0ryt6ub0IhZKoCSyqTGTulZf2
qfCux2fTc/lHVNMpaIXdoGj4ZBUT9KlTI9IB3yIjDWoTlCY0GOo9bTIZMygmCniX
4wWBGKZUjBDwIuYiwtpzgDT2SrthrsbKvNhtZNzNDm5Mu1agzcIIzEGmlcQ3hNd1
qQgHysVbJOOzLimsvZq3/XNoxwyaUSkNkM2OT7FG0ckpP2CtTOe4VfrrZWZyAcdh
pkQSTJ4LYXTjIj1lt2YYQYr1ibx6cNbhGoj4xLvjNN/RdLgqh1LhVq7j/+BxZA9w
FR1G2bvIZNGYzMHk+wIKEynQ8JdUZEvDe1CD7TsQF1/QkobfkG5r5fE2sdf1JjaY
vZYJmlXDx5SZ92hUT6OUfApMpSyp2x6PRxb2e81oGMw45hhfBr2ZVm3Yt6fMe+jz
/mMhQgHrdaZanYXFe3i4jc6AnbAMVIGbXz1WGSSUNxp0xczJEzRdE5kaMnj9OKEB
8xMprzSDWZ4OfoT7kmH0xGSB2FKRZnwSrJOLVx42g6YLL+YUzF9LfjWCoVCmWcEt
c6VTPSYTueY+A+nG7PYY5hc8bSecKBMnhmqCXwaF1sFuTkcw2AEyzY2BsD8/prmD
oWohYkfvuY7fajMLQajy57GzG3YiF41/USAXmrBSQv+pqkt5HxO4XOpEn7X+M8n5
ffhV0cy7qXJeUyNI9h4UacPwrzWUGi7PwGC/a1dq6+QsT1n3UQeMZ95whm6gJYz+
SAv/3yDd2hZpIU1SjA57h5Nfz38zTU7pgsuoCr9XB0ORFUZ66qRKiGTlS9yr//0y
ZIflPcsR9fL4gsMA3O0RiZUX4KKK7Dmo+T5BTqaNntBVGJD7vgoGxg9WmyyX4unA
ze7Dl1Jv+c6IrlQJpG3tFr06w4EWKu5XPcFSf9IWuVtU8nP01e1eBUXtFEM+lLEH
nm6IlfMD9UdUw0bL6c84G0YBDcdj6WQYjabeMUzNvh5CcDU/6IVO+vXqlVb+tCl2
O+v8i8ktg/ezNTa/iMLtztFmgIJvHk4M7mGiLx14BQxcuFgTEWEDOLPYEmyXLHIm
3O/dQG0a7pTbT/d/Uei5z6RJjAJEhsbyFBWJkkVaVgtQVjzHD9NRsoma6CV0Ujtv
bLlTtWSkNALckJpTLZgfkZ0Cct8MXkypBsX/e6miktfg5MwkfXh76HgIIV3SNinv
vK1SIiEolTXmRXQWS3QGSa3Xyq/F6r9ExK2OI5SYe1NXda81w2G61I9RQBpLNAxU
WyzrbA/3azqSPXojzQMomObJh8Uy6uL/bTd8P3wNZkCEDW4Y1XW3ki6uuxw0286V
0IjSyjBLSGOYmAH6rCiaoQio1XA/SR59KBRdLNHhLSuQ79+ReaaithsCwYMwPSoJ
AQpmkR9ItHUXJ7HcY0pUEASkn9W8EvZ7C+vWeT900aiRHJVPf83Y5sDdOFd8fn55
BqodQ6sF/Mo44WfzSSgu/uzwTdO6AUqjecm6EX+ltugkd512iOsW56MZvesWBUAK
fSMLNqy3bxOLba6Y6Gak2CGBMSs85UIXoAda0hW3xlGXoCW/xm3bGUB+//CeQCOd
tnd0EsDmsylFcaOkr7/eJdAgRHIGiPkOQiAhU75ZA6kZnOA5SEOSdUqYcMPUExyl
hxCCCtnERQTt7nCddHpY3yWP6s+/qrTFzfnKutkkAIGwJQ/G0vTJX7WmrsOl6sNy
ZczTfQydTTLBWmZ4Tq5mbTQEgOZhAAwOcZCkO0RNeOPKpwxX9OLh0BJALnZdeqcN
znUVYj9LXzwXTU0mB7ZW3LGe+gvR227ZHM7EK0QiOryPnaffBSHCcrO2d3i6fHRJ
1idAkSGgBAOxL9gdHXabpp2ie7RrXAC4MO6evafUAGFf/XleYLAg1PWAL4iCmOSh
XJoZO26ZRQFv8ATAw4ZEnThZ7JSVAYV7oTXckKIROoDcmF6a49XMunx2HoZcMq5e
pld7uSnH6sCyubQrzuTQkvzcIq4eY9RkFngE+D6ghxOM4nyKi8CajBgpAf2gdD7p
MqXot6LqTGD6umDf8LyF9nqkdIGkx9AHSixut2rMXH+aGEAHauR//N2EwcrUbYnj
hh8I6dDYn5QsB3fVmNhZrHsSPEGdm9JvMAohFnUS3o43Nhweu5EXOdLDzXH7gM0M
N85AJh7GPmSpX5rHpQUvgSF7dF1UmG81few2no2rp9MW9CJegyQhtmmfhH14M2qQ
K05cF+Ws0CADrWNybbeClMqyhsGuWUxgIpbs2Z8f1lKJWkY1SU41Ttw/GOzFConB
9d8KFl46qirqodKiHwLEASuZ7wCDwcfYPTgkUoEehZzlwGq/h0xhUDjLl13SweAw
eKIoT1kusQ9o881PVt8ZokyA1QtXrz2x9azHsoIqNliiwWg5ZXI6/2EPXw1niE2y
hWaSwt75YCCbSA75NWEAoS151i6BzbmlFoo0NWeSOzU1LRbQV3L5Ht6suOhGSAqE
U3UbJcYdYUCHf38+rBQJWdzta477qjtPZBDM2a33gGoAcF0mdAjoO0N8sPjo0Le2
A6PyXXw2ayA26cJvJ4ncxmAAeSTE5xsIaPcNizwxgoEpgFSzmb/ZpnQKPaULvYJl
kylZp1rpkcCV6WXVsh2iE/fxUWUl+oXg6FgpzW3wLnh5ApVMF+nY7LGxY7RL4SN9
Yqjp3WhAZzKHDBszOtUEhy/pI0OrmzXpg3STLPNrLI1hWZeaFrPRL6tPE5/nPLkZ
L5g+TUkSDsXgTQ7kypc0bKu5j6DisWpvy3IktXT/NVTBKa2wSxZgysYcKTlW5jOb
tE7dfz+ReientNBJJ7352gSzGo6ZXQtCOO0spVujcnuDzXm2gKB6KSUh2mknZ6M3
l8kDSrVzxJEoM9+f5HetE8Sehkbkpd8rhb+gb/gmWmrKWxEp1yD98fYr99bhT+Z7
1E/6UoAMvWLP3daCfMfKKx9mdL0aaohhMTYFBpLf1aNeo6E3qIWmSPxAyelzJQJm
rY2AceylIm+z8ww/esRXwjvVtwKXn5z/jidsCLc/XZWi114hxOX2LX0GdWx6HFTw
hz7GMEVx0FHfyHS7i4UmF0OuOHtVjUrZJUVZyIHuBoogLJFZ8IZ5ZOzmuJ/fkb2Q
qkD47CdaRw5aEO+6OYBkWBIHQL4We7q9uqi/nV28jEwPzwLu9nK0NUtkCzBZ3IL4
hn+XC44SAD0qaQDGLk62pzrZ+F6xhr+Nmt5g89qRG/vCVekq6Ni18jRcLCZGxO+G
EJsB8Bj+MsAgBaAKBSV/d2jpfBIVNOMuW05PhYTZe7N2SFcGuPHDTC/A2+eKZZs/
d5eOHTu4pCsHlc6PGGrZJGkn1mik3AHEzuIgEqxPbrZMW8/4u4V2pmjLqyZfwZSU
lii+ORHEMRYRfdrpJ7Ls8u5zf2np0gDHX+QNg8oATpayUjZdjOESlaiLulDt/N2c
Ar2H/Yzirfu5v0qGQyVemltHqNQ1GjKJaehrpjPa/AcVlL61UucegxeYHfvz0D79
Py274EdKuT6NHbtIEOW5bWRno+ifZLroeGk1z61daBGoyauGcxSlGx3H+kqunfW6
Gf4cV7hd6BCtlJDZOZq9SPB5wkdGW4j7Rj3b9qx5zEAzWqouxW+NjHX72wgxexsu
fJ9nkYHFflYWDknwYGwKXZD4Fe7oIhvteAnpHp/M/sXH8VhKrs0NpDIDgpmLo629
nwJiAIyIowDncQO2JP9WboAVyl7eDERHjD62KktaKdDoqZI9YdNJ1wvoougKdN4Q
MkOXZWfwUaGJYQQPOy3YTJJccxlyJ/MWV++DgWzDd7wAH+zT2c5eeWtMyNwagEbp
WL8tKyTLHyLBXvikHAxHLOsbefE3Dk/hgvyRmemx7m6JOLzhT52IqUzQRCswDpbN
EGe+dk4VonTRBqBSHap5GZ81kHgqBo+SD7EQ9ywRjvVFgpRaQYysmmyTY5FHnprf
NTbZ3w8jg9noEPUhCeBz69PylKROfnFPfyTk+XmY57W5oJ2LgOxprbllj2KHyzsl
CIc93sOVH96gZcsQ7TUV3na2uWU+IgdQ7mVxK5CoMKw9kXq6OeE17UY9BPPsc7ED
1oVwEIoCJXGN//IYPoQL4KQu0BmrBJhx2w8Sf2kIo10ZF1iTqyovaYnJJoUiusVL
G7o20RW+HwRH2WjWKxEjJSJRnQMgISQGls0COtQI7C+6LumeO9kSeb+uLO20qwAp
d9GZIqjI4dvP7/0xuuMWWdeeSFRE8Ga5NwvEq3BmTnEdY2yftpy35CEgxEqH7hwt
/1pkn9Be3sQU8NbekuM0vrRg5qOmpw07rhukZt4ya8yIo67oXOa6efyAD8dW5T6B
dkaLdlwhxXKq4N9rfH8OddHmNGc2YNVOH7CL1EYhGNqHOompT4uhXlMZ5nwUtwG7
Pf0aEUV3fytY3DSCRtzUXubFwQZ7ut7Jq2KouslwttDITZ8+goC+Ujd1GzDNyR1l
Hc9Bj3uqBMSwOZGkqTSsTV/GMrfWu53CKOqixNRrKvhrMJtpXeCRysG/TlkCPfqS
sZlYA8YeZNcQBepdwHtWGNXWfRoxW0jj6Xq9rOvqrSJiqqUEAU9jpEFj3uTbNt8Y
OSeGOm7CYQbLzEAd4T89CdgVHpMQ8ewNQ9NE5lSCYkP7mBrlSmdHkCwA6DoEwgs6
p01GyRZSaz0fLjKS5qQuHoF05Js7VctDFfOVAnu0adUVSLBpfbfym8xuCjLuYTUC
k5k5Vljput4KOzWO5hUBttum21Bui97GMobBT8HE1a+EKpKUS5kJGEl/b9BtUkid
g73Ev5vRExxJz5t1lU285EL8wTKql99n/WNXBwgfKrkkz9MDJb+4JzE5pFdZw98u
jNBRu5b9sj8PkvliOwwTCVMnmy1tvnyUC70+K0Dh7lsIdXuxvDKXecUBlgU84og2
ux/4BvWVDNbk6mzljOjbR6U8TG/IiqdVytQ2ZBPpDRCa1L+Jz69QWR+/BETXzDfA
YH9HBWukSJ3jn1959kGCQRM5VUyL77sqe9LRhkVaHR+pf/tORE63c0PyNQZJVN95
6YkuUmsFr1lwGqprFSoZY2xt7J1NsTxIh4zEZLh3yZHYnmujk+X0sIAQMRAzNGvI
V0GeFN5AZb59OAu4V1cv7Rqu7LjmwiRv9BoPDeStHlndYOM7sIKYb/kA4pHrts8d
xXeUvNNpE+BjuQtUI3dz7X0UPd4sTYS255BZAU2nn05kSD5p9PZBoWBU8U5VTDxe
UfY8Gdvv0fAKfI2IyySbyjpX8ZwjmlidGkO4wRgrglBio8zA46M0CnuDdX8zmfI+
yLrUHzkLPtPxIL9FsNEwEk9uA/AFSo7xxp9BRTXFfIzS4WYxdaTEf4YvXve0Yds+
jrNz06VmxrEfkbeHdUo6soAgkKehpdmUfRJpFUvtVnOI7ic+I91Lw0yay2+tqt+Z
lenYbQ+HPQ4CdYAB0IdYkkYmTS008L9PZrqZZcXh08ZtN6fAHKioL93M5gCqmuie
KrHHJIug6rzHuVg2Xm4z8HgczZTBB+AcOR3CXxh3UtjP3ftK5N2uy+FVme1V6qdA
4E3MTiIf1rlV24U0gPum54wQBrNxkQAlhpiUfJg0wwxjc9HrB38hnlKGF7HoJDPS
LWdqM5oTXMlVX/2hFOBLSgoR9ffdKMCiA/Sa6GRt/D1RzVUvLe+GEXr7/T0Jiv43
dzTnTJuuIoA08NA8caOECJfIDa7ZOwUuclbyuvunklpxYRhjxjnn+XS16tziNVwK
+VT4DDfLfsrQ7S7J04kr/BUE8VlL0fkMXnD+F5aQJSRYRy/K8XyB8aP4L4r9WUTI
Vkhfzha2BH9iZqMhlx/8x+jKdoP+cJ7N8WRFQN4F8o8gpSxbXBdEsXW1IhBS967U
yfplKoGjp2UqQuFHQabSqZ4+uGqQzqZ3elLF8IYymx/ZQ3i8tI+AGEp/ZMqUm0rA
zhWk9UY+rMTI/XddC8yhioU6ZY3s6eKjObrlg4cjQUQ3Fvsr5fqgL0bhUSMWhmUt
egE9kkKaKaCZ0XKoqvIqbzW/K3M1QQdedydLvOP6cW7hgJ7MHqPAxcc0bFxQ290o
fTaZEyD9aHkJ2SY4kgmFqEh2dVygw6Q3b/eDrWH561eH1zF1E+H9cB3eiblYuDgZ
wB2a6R99hs13hO8pz7zfEwo4/yYS5/Kv5Dnsg82bM7US+UGHYeMeGAbr5d/O/jEO
nuDStLNHAPQyP2eVnT6C716EXSOO0awcBSTVQkhrL8KO24L1M1Qft27rE5p3psFE
8+mLhYf/HrIYB3E2OivxUQC3ooSx0XOTW/+1YIx2vIQHUIXMPsRFJmryTDqZ1j6u
epc7C0xjbS+jHipYkDZfCCshJBiIPT4n+8QqLVMuNC3sXi9w5ZIv6siZIM0kGB+1
o7sogifnkj6eG4vUolNx0XXykJnTKRafFtfLF8xCTbnoO50s6nkVNnblFFSMBY79
kVG77NGfTQi3VpolMVD4n+cMSsPgB5EWaGub/apB/VHntiV5HyU5q/OvpCpu0or6
kq5A5T6nPknRPiBWKftAKawjyoRBVkeclWod5FmkAZ2snyD9Vx7soie7NOzBv02Q
vSNkTce0NHBnSh9LjkpKzFiQRlh24gY5wXBCDkoMQsniEw07k09AuUUsj8nH0T25
BEFRg7ubFdPzVWFdI2gM8ICmkyKJpT84VJNIhfkgUFVXVcXPWdivGyBXJ1k0SKDw
3W/Zu3j3tsFRLHavbSBNtrAKelsPNY8FMORRUuJ4DxrFNJcS4BqT4W4v8QYIZBGt
aIZm8e68RGPB+f3HZdRerjgG2spKfx3D705994aS+oANPLaHOuEI8XQZZGS3AVUw
rVrrjvpsBdVNX29xSm6vhIamGeJvKqAX0qm3TsqLQQT41jBsDE3uZ55LRbM/mTnm
0G55dRFbBOgfNlh7t9V39RXNqqbKmu+3BFnhA2nwMWh9J858zzuriwgM7N1Z1pvt
2hG0WYXebGwAfQ7zboZ23g==
//pragma protect end_data_block
//pragma protect digest_block
yXxoSxGViT5WTPN2nJswED9hRjw=
//pragma protect end_digest_block
//pragma protect end_protected
