`ifdef RTL
	`include "NN.v"  
`define CYCLE_TIME 50
`endif
`ifdef GATE
	`include "NN_SYN.v"
`define CYCLE_TIME 50
`endif
`ifdef RTL
`define PAT_NUM 2000
`endif
`ifdef GATE
`define PAT_NUM 100
`endif
module PATTERN(
	// Output signals
	clk,
	rst_n,
	in_valid,
	data_x,
	data_h,
	weight_u,
	weight_w,
	weight_v,
	
	// Input signals
	out_valid,
	out
);
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
WNnBs9kUplSfLwXMX9EK6sFI19u2e3pCTEfnPz8zYSe3SWaQ6Wrv+UVMoWEImM2n
HS5hjt4fjs+6udCM4SxY8hHmOQIcJnjfy4/g7pDHAPzGgQm+5AOzpeoGfRybzKcg
IpywJuM43TcfB1rqKsqi9WgMz9CbJIJlH6gYtMFreH52nJ3YWkFUq896Vbz4nmYz
ZycvcaHaV3v9e0lqF8DefEdPUKqSX8f5WlEnWT9XQUl7HMji8/A6L5v4i0q7arsc
gyV/9DZjB4qoKUhienzjH2Uk0wTcfC0wRLVYtf2BORp4BdWN+L+UiDcyVa5sBBcW
hQ9W7rEP+lNPNkTMIG3XkQ==
//pragma protect end_key_block
//pragma protect digest_block
s/HYhf7QmnoBxV6ByvaLmyF+Pq4=
//pragma protect end_digest_block
//pragma protect data_block
mW1HrKsyQ4kCFnGmI7PXJHXAULEKmjG15wcVXj+HLfCw/jHNagNfpjhFjFNeEB53
aRNwNVDHXRClZzFXlI/3yrOrtjNz7NQ6guXdrzEtXgPnxARr/Wnk2rOjwHeUdzpi
Py0ONLHlIcQQz2IUs1s+3v2STQ3X6SI8rg/DcB7JY4dSzMxN4BKbFITXgVOEyfNG
ntzY1E+KvQ/veny0anPCqYaNs+WsXzQPCWQ2R8t5kVqzTcHhg6bHwAFyYGA57ljt
gry9ANAvi6jUXbebm8d6tXPH1r+LbMn0QOJxcrtH/ronoWTiWHE3BLV7EK83pVe5
4LVu4mihTTi5ERk35irm7TM6tokUBt4P/D2LUJvFhbSTimxyjK2gD/e+xSY/pQxB
txU5p4ZpmgR7Jhg9dwS8p8pr+AqeReIb1CUINFLvXMimFI+c7fcEgvbf/GaWdvSz
DAK4Agby4sJ2kJXJLXXcU/F/0Q3FFaXBzn4FmcuELJudxc+76gLh1OqMDTo0sFya
t1BQmHRpf8pq5WoGShUzupPD3UeY/3bEsrmpkdbCTKb87QpR8alrO87dzccls5SL
o21YsK01ApaIKMW0nCl4X0YEWgoekrF6cPNbUsuTHMBJjbOt3QUBsXCAsk7FpDpb
I8DgTjYgbcYA5tqUUrZYKRJyRksMKWiIFhXd6VZmXzI5mcs3xU0H7ci6VMTu47zz
IOtc7GTp4Y514XYdv3bwRo5sXxMEc4fg/VDU4f3GJqdVL1lDgDqVA2MU+/WG2Bzk
JeoQWu457N+AddgW1mDqaG6uC+mkNOAsnTflvttnc2kGglaK3b+nUpKWkSLN5CJz
rQ1oyidMlFKpUeFs3NR0pWFvm9PSWDm2ko/f6kbZcDMEpI4y3w/HEOMU3R5hGTUm
kMORGTsiyzF+FLpPnEujHy2IaQKqlo9yp5QkmFU1IYNql2ehLTOZBmKkYeE5LWol
OWcqA6UpBIoblH/pnrd9LtHKRDnAqbbCg891H0nX0BGnnoy7UK+HaR9n+M92YJhw
QpAMLurdCmqbpkgwXO5FuF5f7DgjpLc7o4STXThVaitrdIVG5MzwHR6JCSEVETtk
dVHvZZqQuvj2mE6JTjXVSrJmkys3MwibcHrN/8TvM2dzJOllHtCPmj5kG8Y/Nppq
6tl+yZmWeh1WTgU7XsqbdjOvYy+gZKtjvo4LDdSrgVETnowGlyGanb9kqFpW1Ff3
EoHFvKh2GlvA1Ti9WhALPRizikoyAvAytEEUDVxKJ09NNWwbjiPDyM4ao/cvNeR2
MLgkBeJBu9gojtN1TREc3X7+v+ghcqG1RPzAoy2tutEVryx5xqbDP7tgpaXkPb+T
o+rwCCVBaLUIru1T0mnj7qq5QXRUD6wz6JEUAtY2MU4aB73nugO5vXyk5orDLBJl
Ua3ax3bnV4sV7txKD2qesN9u9Zio14PryUJc1IPrXqdarVDmi9cI0TJqDb6gNub1
Py4/EtJastIaNiTluA2o1v87Y7T2ZG7di0J8Yy0d6v/AriVRFye0rJBpPdmUW6XX
xQXxBJANBpe0jM0aif8x1TV1oAy2jWbSGyn3TQj1Ri0vwdcQavVewuQkBDaIjeuc
wiZOCr5pfvcKNP21UkaZRjWxgBrlRxwG54vpz1yL8E0jpRObRTP1TlA4VX8tEYeX
keQyc6qTcxytvOvKBW2H07wFfwr9pDmZLCyq0n3nWXnmOgVE3G0PJjCnFXFlcq5P
7O3rTZY7gEc25IAkoHSE2Jt1Flr9PJXNuCZkEj1IrA940YlkIAh6HbQhThE84egW
B/rLvAsI47E+4HiVEbyWNQNWsE6QLENOZFNq3Gpu6RbnYGcZpTy49MUJ4/WYU60s
NVQuluLW3up/zEAxFZPDVBkjnEnalX+2H2eKCHXmaZi0ehim6UAe+HfzUKpxfKkF
vPq3Mh9fcQa1srwRWCyGM3J4FpRTl4lpocRGfawOiEYEVIfXbFrK8nZvGOnT5XKa
AdM8HkFy0wysmoyBN88rE2f5yHWLvRr/MrvUSGBVPg1YkAwLU+Gh3LAH+pkuA/Xx
pY6ZwUzQUEnPYZstG/GumjwCBAvnoagwTav1nABQIv7AMR3BwBe5v1yJ2ErxEHki
p4vizwyWGfBtWiKIiM1gk6AGpSGMWx8Rj4/uRPoIssVaMCZkRLZwrYlJJVs6EEZF
mQ1BfUQsetdG+M0hZKScBLUyHboKqlaZFVQ5NkRM0nuw4H1Xt13sJFY/7NgoVwkM
FvmhnJSyXys7O8Te/KQw7zryAB2z57uDz3w+bvYvHCnxx8LdEDwrE8iI/YUIwiBc
mCr38tXZQIqKA/G3WveQ8k5IswPWfX0yKEJtQzSX7I5HTAtLZWekegozHd4Dmks2
5mbebtC8fntTLSXqds/CBQjNhrKrc2anhd9IpAuCAoKWlCZxmUvgkbfjQYJbVg9F
f5/s7TG1McG+oko3e0qrUvL5+R8/+4GF7XGFUdnvtcjQ9WdB9u2lnbOxcDm/haKV
9SxTXqHVzEZCljZetEFHmoHY1r+EZQQYBhss5Y88cA633yTrnVdnOtp5KYrGj/b1
pFd7d3xJLVwJ9rZHOGvkGDr+gw2FQGbmF59ERMRN0km+YoBgDL7p5lr2ZjIVkv8A
NpytsYC6n8filHxX69nzjkPN64vG4t/5m9uvtZg2MwDYUfkWuAntD2v3eHYmwudh
v9eY2pkzfka9jjER/HdbO1X6T0+M8O+LJhcjBnhg9O1p5xqyCirI07EA6wUNhrRS
F79+7UomOlrI1o+5z6x5xcsxtOkoLYFwubdhSEXez/PXeb2g0qRTDzlWODkLrEZ7
SW0aBISqO7HC4ZbEzHzeZtKtOcIgEVbmUJUpHI6E5GssuwLyG//YkRSUe/Fi9+R0
/qzej5I+F1JY7qsmufFtoH3en5BJybhhwTbPKtJI0Hm3TF95E1OCZ19REA42sRpo
JoPpD4zH5hxqcRmtPJjGkcYOt7jFQlCiA4yTcnKBN9DcnjOnlVgqgEAnoMUwZ2zN
t59Y6R4zliMZicB7eW++kvWaOI2r1nlBb5LQ/byBaFwyjACRG6Q3HOZchqEroPqm
WzbXXozVSRlNOBmdMcKjQK3mS6G4BJSYC02xQVpmf+Odghu1+ACQpFouGo7yB9DW
6Aub70kTDhI9ZhlZPl+hpXU/3Q+P86l9Tld1j27s93LKVE4a/Jym0ce0QUirIc3r
FKAAME3ZnHL8nz2DdbIgIwssSqMfeL0XV6Obi68Ie7N7ZUvHwuUgFv+E9eJZFGkH
zEZ3vdF2c6ApaAm31NNlUmnfY+VKIyLwtDOp6OxNwaebqZUHShPuwqOWLckUCW32
KUnwjfKo9JM3ey4yf2s8Sb0OR8oL09GXxhxK0tIVoAWO5wTvpI0zNpw/vrv5HpvF
A91PCQNFeGvh7MVjWSk+4OJyYRP9vF4aoPJZVPns/AgdYLZELaW65CnOPgbXDmLT
YP4+PSiuGTAF2vhtp03pfuyu4V8Jt0IRGWrd5KE53ji+39aYN3JVzT9HVV/XFkFW
GJk6szGRW6ulskzIgwcYZawu67ff9pTYGHxx4JLFKxYsRunkD4YLYc2DI825vMsT
t75Wjcb1KTGSc7b9rzbTWLiIAZlTR/aUmTfBujxAU4n8S+/CSb2pGhgcd6YB5Xct
jPYwssM5ATR4PV60UbpJ0VmfWTksgoeUaGLvdBgWsumTYLaaYPfGa55Q95L+1oz7
lYNEK19lwwvwWjm8217L7dv6YfTClZN8wGepHFRbqzO5O2BXRi8NHK3346a1WrL5
mubXgfaBB8FRzEdBWvSNca7NG6awUJ9JZxxivxQ2iYL72i9MwsgBDwlLU7KM9Erd
vMiTiVmy1ywHXGRm99WN/iQjMlAzreSv4PcMEU/4tcbEVWfDj3lmUQu4+DezzCJV
vdD0XDG7lpo9XFLf1QkEL4DkTVJi81CyQ1ebJ7j3kHkObfxB5n0u2jOPaDA+l7M1
8ZtA8j/S9d3DyK1Dcr4xubG1YpYXByJMKdGdF5WFXuA5gmHp5Qm4Hd48aCzjazKy
6lerMKzhKtBN9xkb+rOLRG7l5j8hJkuGSOfyKAKvPRV4Y3l0BWTzW7wIwsVYU1p8
1EgdTSDaKmNUCd13zf5fHBJAqiXhbi3uFs2nRfACXx2QSY99K3ZGR2DaRQo0lqaJ
NpBJ+LHPNVIVjoYegHtub07IVIkXb1yZMbPA5lGmXQ7MqQOa4oAYb4Aty5BJ9EP/
4ifz2YM4raen502WmT4W1KsuGBor9sccM01N44OujW7wexTXKmZNsYcYXQzXHUxe
XdazHdPsZTtxUl3KQLjTk8qduHDzMrp3yeqTs38pMxGkUUdUTNBqn1VDkNcpR/WP
A9ByNq3YBTBh1VWrFcgv+R8VHzIqxUbQV2a7X9CTo1YWGMfCBAzLkWKxAozI829w
37YEdGZJn0tQLaXPgVcN++RUwwlMVk0/H9bnGs4vyZDCMYLjotbcBwTbvH9GFAVV
e+hnSrHm7ULO49f0Gme/EGK3JpQOx8ACdc9FLm1Sn4u4sakWt/IfEGRJkh7T+kJ4
zd0EvEmA08HQn0S7e3kCevvgvFgQgIE2QQO8LRwRd2MA3iYp81P6idwlV+BZz4/m
pscGBVi7anLzswIJWSWekBDOP86hx0EaOCXNBPKqrTg1pKDuD4awwE851oGLuAXi
G4oXivx3/V4lV9nRcXzGE2Bhj+aSfHzHAQSBqxLsz8JzUnmfno279WtBGg4Kv/bN
yrW0nLsnhv2No2uZYXa2q7KF3X4tctMGtA/uqXaPjkkozXrW5szvFYvcXg935pJi
Fsu4cxG8PwSpfmpO2YEzJU+aAP9DTpTPmWJV2rnXuB6ZgjrYa4MRjMfEwCAEw0ES
6V+k1YQKmaPwbHx0nkCaEJ14JIw88Z4/pNO88AIowKPcYmwdBxW9LLI8tj/fjOd2
Lxr2m8PVeUe2JfUmotE2cyPBiUGuXNx2brLCnBAXM7dtI+5yOHKizDjjnhSHm4CP
JUu0jaeJpyHItJ4uttxNyyQTj9vhsiOBdI/LCLdni7wxDkMX4DyNddACAxQ3+9Wt
J3m50xIuAimaY8w3ki3LsnTF8ioaQqCJmAp9+hSXfRkyQNw/SSbja8V8IlfdDkvk
/9Tte656rQiD6QHUoF0/X6NtalEr1uz/ziv7Omht9iEXBbfKy5rFMV38RHljriKW
e0IfIzvjYEMgOb14sNXXuOQJiNbrkOHePJvI2PqmU+Lz+K3GtuK2POi4EFXb00Fl
Otp0Qh3eoAwxyGrDBwFpUXgEi81lwb0cFq1Xeb3ZkacjTIguGrSg3gXW3dSOF/y8
xuOSe2yF5swlCcLK33eMDhoXpFzCLEQGoHvddJvLffUfTTzh/dcDpUi5lpGKpdpO
sbgbR1+PAipPRKaHMPz97C7KblR/Ky93/3Re7+qTFMhPNYjwz+NYpm4B7C+y+3AY
5tz4EH6bMAeGSnkkxfe9ejMEuzIIenmBkB80HBjRwwqdA9OT0WCoUl8MOEcDgrAy
WLDPRDUwOJdhyO+sOS9VPDhkqxGQMFzWDT7f46WJEpYVSavCMvDdxcjD/jDSlxOa
5Esm3MGSnctiZTC8M/5JsOhE/hjCTiICiMnpgQNul9mkmCv8Q3CrBnsckiIkOC+1
sR1+wd9eSTi/H18e+SMK2PYK0CAq6zRs7ZqdiZPxxH64sy/tDTxpMjkecY/qX3+T
8RFb4bl7xa7OnTfg9dQSP80XoKqKAbY2wM6gC0GqYBlY9G1nJDJGZrc0YzyrU2a5
0+zAzP9VImGdO7L7oBr/UdNZ7J5qT/Ew0XvqqaxavWD9Zjp3VAiMwxRh/GlSTyZh
bhxOYMZx1FGEXAz+xOvvJmoDOOs9hkgarIcUgXLJ2UyiHzlZCpvZOk16H7+uN8tt
h958hXke9Rc8452k53X0uV1H/W6EDbXXuratvoGJCP+6o6X7A6X3bbjRPb7pSrxa
QBeLDJnL+QBmxFdX7S1R4dYBukmDoICiagxqZU08df0YGY7PIs0+d1Rh1TC4Mbun
b5ur1O7LIUjyW7UJ+3B4tyIfl+JVJhhq0d8S33hMtc7NrYgd39s8KFGem7m+Q7xb
18B4H7XEkonMF9ldmCMjeM5gjbJwWWcUYL2MS0yR/LnjAW8tsNqrJGJXIyz2nPco
44aFHQ1E6eMyUtRb/2IGj2Qs7KZ0gbFwrO1JBMmYxQDUu3cwT9F5MOczDl7IKTYP
hQZoHX1JXLjNjuOJWc33i+QZJBblDC7pe+UwSmqR6kPg/tAwMmA/4c+UH7ye0/Rt
ypml0wX23OlTb4XvRaZfMOmbDDVVJ/nyfAhhn+CwaLpCzqipb9Eo3MvAeoyzSMNv
WeE304Ucamt60mD/DWFDqT9LR1mMVry15H6EySMAX7C8Ow/9A3ZFKs+AlIlj+UbL
GoJi/t9D2FNJm9J1iQc24nUIt8DyKyLHfurJiTW+ZcJnKYBFWEBxwBudg9zjCT3b
NC8HfvR5eIGL8a60CJ58++tD5EysawqYE775jFd7j4ilyWJ3sm7d6PglnCogA79h
ZcArFjEK7aeA8J1NWhpojUC0/DiPt5lm+YaCGvvnnBBnWa6XDIT22cgNvV/c88fl
Gcp1zuQO1vPEtnjdarG5INypZtugNUHVZkgS/Q5aP/nEU21MwdrriJPu3BeHomCT
QjQwmZGv7moNssRPHPKEtCLrKO5fCWhveJ44uSTgqsA3W+SnBe47iwNdCwOrDPmV
plLHhEyuplBbCwADpnIZQ4ktPAfVegkK5Rm0liSZ9S6M6Mfd2P0ikvULejH8kZif
LxMuw0okMMeK+oYdvGCAFCd561ucN9MzEb8ER3dvoJqZaf3jv9OxeSE/IyVJcyGf
wPB+c8i0LuY9e50Rd7Cau/z0uq9gPGferN/OxW0TD8CQDCCbrjeu8+xhbmZaA8vR
TuyJdgkwyPmmrrG9l6DCkH/VFzDMzYIOxxzmmAp0Tl0B4yMGVb09nGO++XBchLe4
/lHUZBzQsAmvFDhBKFfjvVxtcLXmfCjHv+BO7bNm7mKZTMcyz1JApQFZqZDAQD8o
W9gEE6QA0wl2Jr9CLi0N4fuydXBki47u3EjNbTUHHsyAvSOjVuAt4erapKcA/GDI
PgjtDtmFl9XQ2FhbfqkP/Dy5I+a5TQs7FgNfWEHjtaWRBjNgPiewNBKgvhTcZJy9
kqchKB4v1zi/YDNcAfdlASpAyofZlX25LZtpHUrK+ethcI6O2cOqaMbBs9D6TpEK
AZio8qOO2CrJ4I/PRyes8STLvBGxRBqrVR6I9Nd/1al9slI1aa3H4zMgL9a3YiOD
7WcggGvXo4YCfJRrsdWNz80lWRQmdJTXaJcIGpVf9/UxXCBud87mmtGS94wc5US/
jhOlP7ds/koW+gIO9oe1JI8iAHefAAwcxMHMlJUeGLgx5a8LFp6bTCxhN0cMsYND
4Ox9LtJrUZYPL8g/FEQM35P+ldP+KvobaomusQ+e0m6ZIAYgFwCX1GbdTFlPCLRD
p8krajKGjb7Ehx30f+XRAiItV+1f7Lt4XOzLbg92IV11ZADQNrF9Wqnf1ALUjpdZ
9cZJRW+Pv0Kp9ZCncEI3vom600e1pxLj7IHy43/7B/t2o24tFFOPx8LNjWcsZjlQ
o1+O+WMM1Cs6g7GLG9p/Jz11rnFWJgAhdxqdcox/h205aPhQucvAEaK5Zf0WkCZw
51RFxSqf/R4bvUjPLMQTTEt97mwbfZqCyhwpu9AyAQlfCM6eick5HEJNH2axApLY
0/7wC/qJg/GCaF4JVLBNHdAZ9q9h3RjCOtC+odWqBvllpvX1Tt1Uu7NrUsRBr787
GqTLuyV81uNAhvw+3o/xJMIfFeVZxrGAO+DE5XdXnBvZQV97xJHcPJhdZL/efXfY
LezksCv8VGPNt9GZQLcXcAj+dDH4BoD24opmO7qvaoGaY0HtD4EqY+CgQC7EV0dI
tWNgMU48xXEpKERNvBqMPfZr29ERIG1vixEKN5C6DzjTOWTkAZw9qH/OIoRY5cLp
BJh331ed/M1yMKZnWjBFosKUoo4h899W5v7byuR5ml9caV5bcmn8wZf9h6ipGRpe
XQ/ZMavixECY54PbMqJLFd8BfA7Lb3QVMZB+bSua11E1aVj2Mdjyc5jIW5TiJ10U
oGYx8S1j+POfmH8fVbZ2MbBxplQtxbeP7QkuLea2ypCOx/iJpPzNmfT3xyfv7Yc5
hechbUrq55FfEgZlc8/2Lfp1Agkwwf2IjleFPY3eo8/iPgMlevQ6k8Ge/9oyxfME
vGIELTa0WATGhmYnotxlAHQ1NPxpT9RNzkh4sSnfsyK+OJ8Ri9v6WytnGrpm/8rL
VCFveZ+YtQt+JbZufMlKHpuNt+p/7z8WInVXOFr2L5CLej9c5iMaxGIRKGZ+OSVT
Gzp2ofhvCKrXYDLM+8yaTBw5k0vnbnqPFZgzY507l+JcPcN2am6Nu8I6K1RAi91q
a/BNOegnI0lfuSiTJGtd8A8WQBOWqXWuRxTJjENYueH7eEtg4fnB2zgWyCflYHi5
k8g1T0RxUQzwWJlHJu92qTXiXSchfC/ObjOSaazmDoPVFCIcFkqKnUIY9f12J9cK
jcZLBQcVDmpDTuplgNedN5xWUT3MWCGxl10jYzFE9rPmBgmgvW6+/vgAxhu5UZxN
/lto4G9vhFp5bnfByWl8Jo/+UeDqTx3mevBNWejnYWJnOpSp0jN7zHRc9Gjxf/JS
RnHbcpXedZEzo2gFLIDrvoru98S5uNmdEnZG644AThC/8uwI2doZWtc0Aoivyv+w
o7nQeb0YDRKF+xkZmpRPK/aGEwXvfPzvNdN2ooxVJTrtJtigPNewn8f+KEHVLRhC
yN1qLmeCN+SnbMFAfDnCqTiQCrhImf8+UFCwk94KLmJkHRGOb4FqKwPEwbfovuER
w/rvThurmZHmRYZ4mUl6QyzJ0WdPO0NiZytjnnUjWQQKgP5rJXJRa9OmwCiP62VY
QWwZhtQQgSZ4MbcSwiKwJooNdg7CCkKNdUdpvo47GmijAHXW7SEeLlB7q9RsCfV3
S9Xn/R/Mfdszg3bsb1C3VXH6X9KpJmYmXhARzipvizTolAeXUNsJgJk1hxdy6nDf
Z0YQkPWk67E1myBYOpjLKbvcDnaQU4bUzCDpnPhWUIwKDydr5kOxMsiNdVVEj3ak
xMVyr55JtdWpjFedXPqRM7fq7ZAna4SjtZSO/wkG6os4PDDmu4na2JCyMywNE3j1
pqx5cyBfNW7Rm8xeig6sXiB4DVjnVm1VFh0Re/wDm/JwWHxasVb6ndH/vi2V4Koy
GogQO3qhxsHfamnAZplcK4N+FelWCtwtoPPL0cUj9tI9//sD3VrfsRtRt8h4VYf7
50b/aZ7P4v4QhmRDKX7QZqbOKuxY3wfZ7VCUpC+ckc8HLBtWPmQAMN46S5ImSMHQ
NnBK7cR0cVm1SnIuEpsPWuYU1b7d9C9GutQuVueB8gF9FYyvr5Rda4FlhA4UNWYL
NzqcjzF3hAPwPML9/FH8xmpgVU+hhLojJuoO1uHU9MQH1Gb+k7jyDaSe1WqGLD7t
PfSwKCP4eVbK1io3kq9LgZb3smiE2J49ehO5D5rN9dBI/1eFE6/zoyZPyGWCoGlA
K6mL9wScAAoBxmrnaFkfoGRhPDn65pXOIVSyfXkB9bE1N/QbEmbMNKtDgrSplhhS
rEW6VGWV5yNZ51181NTgbdTFICYFTUPJPwySXEXYyv8bdE5n+oQciLK+una/dVhm
2yzf/o3I6cybm81WCcE+Xn4gcwhiIdh+epFusZHMcJFJRa+VvciwcUzJ36ZceDx/
iHawGUKrH9SLkxkLNfsqgbn/zWNJJf5lGYkZj1WIALapGdBS+h4ZiAhZvA8CHev8
oEbq5/fLuFzww4tdlVxNnyeIAyYrJxfwtq/wZ6WXqdoCWjmT0czOw9YTsSoZL4gh
NCI9IC5USpK9bdOEUmlkTz1OhwC1nJbnklNpCK5KpEwy3ULjuu8UEVvdZXjJLuf5
ZIH0pVbJfBfhDeLEsgyLTzZt9YuGlH95Mhx27Gl3OaHc2dTAG/TTs9NZaR/c1p+R
WcP1EbvqsApEt6yooQ0WVAq/1Dq4FdfV7DGoLFae6HWXav+k4WmBRixUXp4O2zML
FOESKC0Y4Ym13kVoK73cMaF3bjyivzOgD9307VUUrknhY/kgFR5eF6JgNLIobveo
aD4T10Nb+O8Kqi3cn+lne5wWJOTOmbowoI1Vt353t/VlqbL5qxxsZEz/jb8YrZNz
OmT+nRhFlVqbqQDhIJYJDEmS+u2laevjwgfR+v4gCI7ZdmnK/y5a0L58FJJ5TccK
ouE72IFqy2ASAme4+yQ8LF0lenHU9/hOm/ZcthdPLaGR40eRrwOtd0e4OnGl2bf8
HQsJ2OPKybYXm9eGcRDviyQlttjb8TJ026LZMqnqN9pxZ8fGjTK62t9k8JE+7hY4
VoeQdWkVG/NuJoEbjbVnVT6rwszN9zsS5asE7+tBbUTiXKUi1mS4a8qd90oNfHBs
r1EEL2NKeFyYkDWPkqNy/FQjjyUY0iDqsnt+QNeHCIMI30x26yMBLMeMdp7A644M
nVIuNlA+2M858n7oL7CAGnHT6RElJxCv3joUGMucUVOnUzDlsPyNJ7vHJShFRhws
AGEYlTRMu21vBfq89iGeET9X0w99x2+e4rGtY8zirQOwVL+MSaykSZ+IjpXSDT1c
FqJcsFdWg8iNtdl6XJeiuy9gS8SkQ7b6xhMS1Yyuzfd3Emj0/ufJsskHYvk+ERw8
P7DiQCzIqhDclumTKAlgZbL4UfTbColowe7BzX6bmbIPja3YrCKewVI03EOiahdK
sxUR1Kjm+IEkS0/H3avwvTjW/M8PX80gUIBA8PM+kLfPnlwfCD6voAMvKoYxTL4/
I5iOGw7Zxy89HylBoUA8/sB7uF67swca7Ur867GrDxT0l6nE68pDQCgpDvhh4BVZ
eLFqeQYpuamQNhpR4xlYnz8F8HwYuDaGkA48/b/u0xvCDIGo/fh5tyx3cmLveUJh
rBdWlBWXI/lGYlNGOZlHrNbVseZjaI1Dby32yGnBLoQH/ywG7ceoHbfbv03sK6Zp
V5Z5Gh78dK8tas3oxqzaSzlCuasbMdeu3hWEY8XKzevbSDVEC+urFoFyxd5KX33E
E8gqm0v50FFRl9Hm4Z5LjXT6nRwG5M0sMLbyl1cHJq8SNfXSARdp93A/A62u8Bld
cXScmiQ7giabpkiJWT7yTgsKkmPVz8P0gfsqh6q2078MYYbaEkQc0wYGjLCnzw9G
8Lae0hsdS8cA3EPWvqcqmXHz+iLL6O96OcmKvJFXWf5EkhFAOGpJgtquTPDazAe+
eZE0SaWFxl/VkC6gtzErwNp90uBuwoYxIRRzsb796rm/4SFnWV02gdiTGpG0ltZ9
urJmZe3/yu5tqBJBTJ3zxDoR+m39C3HqQxZTK2V5YYCiRr8oW/6jFj7A4eKgefnG
NFTsOS0BvdiIlLML4cRArqKCn9hr/BED9RyZRrSX8ips8u5Bbt29qtDcKo6pIoqN
RQKNIfDODdODCuTDApazN1BvBvFvM1smrFg3f7HGFJkGqAcrlZjtPgesgUl3VP8E
o2M14iVkCJp4SsWa0SkIsf1GNMRTfnD26dKHdYYgZZ+JEdRo/vzjuHctUxGu542h
SykRikObucSh9qNGdyNmf17pUYlYk6eaBWXFTddD4LmkIegMqwnvfZUULSAwXXKb
gPy8AaD9BXhml4+eiALPc1Pv77x7wZv2OPR8Edua214anT2iUCJIKqY1bOnCiHcz
Dh2d/xeE9F18lWko8LtgwpX/EiIen8gjyvDOnAnx166og23hOWmB+I5unFCzxHX7
dzzgGHmCgqjMa5fSnfcE8Xf6ULHKk4nFe/R5yDwb6/HDaynRx5Y6I9aRIz/TKG2r
9zIEczFtVpXtIg6ghMi7zzwAJoBHZxj5olcDxwIbZIfOG5vfb/UOUjU8U1mBu8cs
vodGm1OwdZbTrdVpvBJBKu69kYdPEXGa8D7qujrJ4+7CvMmLuRSa34aFH4KdaAg6
gyZ/60qEZx1phoNbGIAEu/a3HboMgixlhvJlXyDQeYysltKsaHofTI6FnVsUZPwc
Kc1w/hF6WOOuvJUFg2tt3pfCf58YxoNhh/UwZMr4zxBc5Mt/aQJu9qPXhqy66DYN
GSDGTpgj39LSkjnWHeeXuB7UA51NolEu03zSHe2AMjduBWyYIpP3ib5NQwtS/kQr
pq5SVE64sj7PKjVI6n1f3bXbwIGOEU5hn2DLT4bFhj09YOUYE9MMP6eYEIMLC/u4
NZRd4pEEuJBfyGezqcHtpgKkM++1zR5YHjT5bA+y23Hzk20glZnyGUPutGZ7ebGv
vZF2YSwjODmHh8RmqycV6lTwCb+iEcmmYO4LcRs5u97p8VGpK3J6ZTseEBtM09VM
AAvrDQ2pC/sJSQbO2WrfYI5+l00URp4yLs6n0PfpZaGYYAw/b0PbJH5pvY1TF2ed
wu766P4QeIQDYRv/qwsp/pyhE/taLkt5pHdiD8O/wO87H5+L0vrGhCbVLx5ghTPC
X4Aly1SylYPRdEqhfEyFhrAJ4aYZiDPy+a1L6t767Z+wHRtEXdzZcnCQgl8b2eSm
5xgpRwf8TD8MKHnWFIkfOWlYSa6aX1FU20KiO6uAqNtgR/fxEQ7bx97gBJttZ9Ix
SYTGLPaRVGfZoX8O/DQ0UJYHNC2ilHcXDOYio5LksTZbLPgeACXGgNFbdAfvZocO
LZmsQqISCNseFvWJdNG3l2tDmakpGP4AdZZq3ct/ssU5HwFqqCZALpp+e0JSWvBS
Y5K0Y9J71u3S80GL2/SLAxXDMO0mEN8uH/tMfkmt567UcLw/PN6uhWqrXyVornYZ
jinIE51376dqhqoHGfTakF7sMIsMR+8Mq8q10cUic2wEkAcsKImoRTOqMeGyBPfh
whenDEboBUTWlhdpPDnprtIM67khfcPwhH9NIudtiOZ5eVh4SZHY0DzPYT/xXRtO
WbQVZ9nooeHgm+swdExuzjV/enWmqeVuaTsbwfXpZ2yU9vvirhNp/zk6qVkl45Bf
Xm5iz7rSg8eExJ5se1uAsm4MlWBywdzttSXk7HN5Ia+kbxTIdy+I8vexIV7gQ4mm
dZoAtX490SoNwwLwMHqYEKWpg2V/aWH7NQVAYI3/vYNsJ3DsPFU+8nSrlOlOhxR6
xcH7gOfGhHH8TSRMClaGHW0qg78aSCvhhOCxy49DGqg2daarC49XP+H1NQyifU+q
HZq5H2O1wRl2wAPraOCSZ8O8QOzYA8K/YInWbvafJcC38YzF4JexEzIn8aI+ZbOn
A2V1Tldueh8OonoPQbzwIApmCA+Xxh4MBQoycNsppaFC5szukQwyZEOuszcWEMmB
09farp9R3RBiyQ0kRSmGFBRybVTTbjaNwpgIdKuB8TrpcZYW2iyaQ4HnoZUejFS1
MXneObo256j8ZUnnAtVBduKfDo2+do98uvvNPLONxeKHDP/WxKaGfHh6Ans42etR
DeNpOPrEFTosqzExa47aA7JXmi+7rzcJR2CdP7qTwo4SVqPmzm1Js7Y7rZXH33U3
tuQ9W9pXkMHo+BbNQta+lhic3lUVC6TBLV8J41Y3ocLsgmx0Ccyvk9pX/WHJZCZe
PClPzQ8LgkJT7iQq7lb+K5ZzkEY+l8qD/jaRgE7kO2EH4lkzh1BbdIDhKkW+japV
qkaSd0YA7B7E+9pErKSTR7Wl+X8slFwK/pRlI4JzkSkPf44LmCewZZUtPznRhrHT
h9g5NsNu2tFhnA2l3YVRJe2dPbpk9Llip6lJvoyvSDkfhX4fDYAz7xyVxJE85Iy7
rtNxEPuEzgo3/su0HMHCqzo8clpGiTLzK6UXRD+lhaWvD1K+dmN6fLhzs9feIMkO
JUUHnyt2f0zOr0fULrixEoOrrowoyxOeu+/PH8fD4Cc7p31oTS/5Xf90V+87MBED
CPyAC6WXsWobep3rPkoR8EQ6Oi0rYUtL0+4BlGeRnpSQyRvxQkPikNs9t37/rKJN
Ydy6iI+Y1l1WWQjiEW8Q8z6V5kp7npDOhXsWigPRg1qfYKsHxCaaDsbPiiZOj5MK
T1R5H1LibDxoFkOdoW2/jxxtyhuktsXM36uUNiOmIfrvAWPop5xopm5qgZZGL0Zs
LdppwcNtPV/ZV5KEGYOq+jg3DHUMsZ3ZgFhUKylu3/SaY2r2SBW0HRmhVSD9+eXp
Ua+nc4lKQSnNGT8QmY7H3dMLM6luOWr5D4Fj2VSoe0IQcgOGwnUUiY0/xOy5MUAq
YH/tJsYKYrt/yZAFCeoYalGB01fYxAqHbs8kQXvrvXO7w6tO7T6akrdK7GPvxG2x
FuZFfrSSZiM3ekE3GEqOMPlS2hqaIm9VyxqQSBfD4IIeW+WC73yk3cEQaXtloxoO
JwE84eUI+WgBoKS0+nP8ABsen/q1b77WGX85Hsrob884DHxu8vZZ5Dd1zREH5tuT
0TjfeRzUuxisDk7AyjzBkoL99A/oulG1FdEzRhhsp6IipXa9VjlyU6IA7LXobyPL
YTky8rKDeuTONKg23ynuRjwTiI2ZF8W7tZruTh6c0QAJ7jF+yWUc3xS5SILmDNhA
oPENPvB/AooJ62BVY4F/FN/3UNdCZYNBkru9egmASwcVCFHZsfsHlaMRiV39NPGP
QhDfmpB+v836SLH16zqgTxJE8VqyRG4/v+5Scqh/Gy7M1ZT139xjmk3/tRBG3jtA
7lZuUK/cfPfb9XvtAn/E6fCgDkSmIl/klwwlPOaFQawYu3wb9KcNbLR+40NQcze+
kIBFkam9sVaxRP7ezgq8w+SLQWb+5l89+L+L13V5/rhzVkBS41tGoAYwtxyuYACK
iW3hgBcaz4cLvlKU5BSkp+jqrxmVobiUI2zuW9q7C0OEOwcTmqMK0u5M31qQqDjq
0M4rHDqeeJvqlGizPcasLGaToND81M1X64f98PCHXAPnx9c7jAPXZMGMLR8e8mSa
thGEzrZyRRwJqYUtZfWOL9S0FRG1bROzcXe8zA8h6Jk9rkTLIx3qUnxxks5AIiaT
dOD995fWHmy38Q5fYmAEahHcx30QDHIhetnaNlqn/oZE1EoKhBhKAamc43ErNuNh
r6Mruxwv3OaQ/VpgcW9wBwNZIOm4G1891GJ/of2yC2iM/b7ZdtQ2pdM5HTe+ZMgX
GZ5T/c7ayFe8nnNHQ+ZhkMAiyqBGSaqhrbjO3l9YOITzxRKKZtIxDfBSE2EaVJ/B
IhY9IpVbF0tH2YK7mMERzseF1Eyd5UA4rLcNpOnDgbQVhVGj32TZzKdMzTrtULj7
cXdGRJ7evu5ekUDLhWCWbBlMkHdNTDkeQap+B2O3lpQR/vImhQ+dJX4+WlBwjLsD
TG6ru5AlxPveGAtxJSFUSv68r1rDK7X7BNfx7TMCowocdZwF/JWDcJHK9iz7BcY1
NtcLpQZZoiXuNOptznA2D7t/SxmSgK5yPvliX2CObWQuyd6EC/s358BgB6LYihzC
eiUGA9EDUGza/0Xbb3f0cP63PSpCHtjdiyphiHUrKHkm5ScsmBZJNNnCaSgwnbgd
RDK0VKSJymH1YrVwr5Yu3im3aTPAt99Gg80TNCvOU6fDhhO6G10N2ROs1eMqehwM
JYaBPq/9QM3Fs79+tJvjyV/30rUfCq5iYqJap8SFGuOP2SWibMa5ZF7KRtHJk806
BJ8pQ1r/69kUlt5Kw9C2jwy34nMSCSfNZqP2jVXcsu/FukBmTDKcWNX6Ik2WAmVM
giwJ5W+Q7aP4jaMZr3bQvip0m1f29mkoZYsy1QhER1reLKN8GTdbIypG+c0gJQzo
yd0BMYLvCesT2UbpajlYXmHBFK0VvFDEbBtB6VqqPy6U6DZNJIl/QyMULXV1V7c5
h5g6DxIDw9l+yc2A+aBcaTIiWQKOw93iw8ObJCp7WTXgDGKqxdIJpWVrDoLXi1zX
pGWGKbtfP6lpIEWwAwq2ipOvuFLrPHmQOv2915F5PmII5qK5VU1TyYs+Czxwj8dB
MgfEC8sCqmHAisWzDueEqLXtZ4xWH8cK0pkPz+rhfCYFBQchDoqb8MX1SE6/Q6DS
I5xJxvha/XVSjqF+pkJ0WnPt+jpednlVaWo0PK+VB+e1F9ijPL+/vE+fEgd2xasL
pSp/sN9DJSGUAB350XSQ+PbPkEpY9tHJmwf8e4otwhNl8MLZTPaWSdcQ6MBhNh7P
gyDXlbySTAIKciFojpGIrv+TeN4nU869n+hjrr1jRHltVIbQpijf6/2LK4sib8Dh
n5lOHLnHvPfpy5cgxnKtNKbcqeiOdzZ6w8PgTphIt3NvGELRFptECe797Z8B2GKN
4IZk2CCe/DlwGl5kp+/y3jSjmXzUM/s+K56kSwu9YiGxqRfrLnkpLMXQV1qOZ/jP
vZmvKXSKx8137IVtzaAIggL5U2MXfD1ILT+8QU+WMgG2p2bhtSWuzb9A9r+Rkw2Q
YqacoiRjO2tX5GRzsW5yEya7binEyrca/BGvpi5RH/mg+sei6uuV/Noumr9xShi0
cxDBw+ZscVo8b4X5OXhgdNYBxGMWuuyf2nCR4w2IYdpC0OHCL1G4pwWXQp1Sft18
uASuyZ2h9mw4bWda66cXrYSshu6feMtdboFEljCsUR6oXr43aX+ZFeJ88IwfBorw
cD0XJREQBNGB1BHQU7o/afBexfxP4GTLR75WJurw7ViI85kJxgSR+a7jphDHttXD
9KtNs9Fx5nVOZEojTYPsJyE8u+koNKnonbcm3xZpwIa4eEQuD+c4GTaL6WgYCaFG
7YgXEzP2AwApxjWABzOW3HXx1r5Jf7BKu5MJm/k+gfz6lMShjqp48AdEhwv/AZgw
6TPf+rQgKUKdEK5ftCLv6ZegnhSLYHNWN8KpuOtrSwKIk+6KbKrPxeIjprr7OcXV
F5StT1bimLleQoSTb9912EqFFan8x78WKi3iZqp9Q9B8WDz+3A5kir7n2Li3B6dX
OG5lfVERr1Cc+iZJy7k0TcmN+x4nrEiVY2001XG9kPQ4hVEZdUcAeaTvO9qzCYxK
W14CGmuhLdc+twDihY+vPIWt/UuNlgN89aUetDGQKw51vaZFzLoR9v+Dd6CJiGPD
NgcFd4oiGi3BBZYlEak9mopv/5YkHDWR7u2YBwh6hgAsGgZIqQWDnWREZGOjBorR
Cq0vwGz6l+iVS7oWVUj7lI3Wy2h7olKircfVTnOOP0gdPi6FCRadiKh9r8VgOXzF
rKwNEVgfsLmdP6FAnk2SbjD5rcFZrZtzBSgBGAZ77Dbm61UbzTkCV7HD4uZ7nEke
KUmdoepQ7mgH+VS9fnNd2eY8tHdoytZztqcWtUdCZGc+955zYJdSZoLEfCg6cHCJ
wVNByzS+NSQ1R9KdbKf4vfu/RpxW2AUMaCz2l8svwTOR1ajtmR69cQwo77wZvAkZ
KTNSmCVcSRHp4MJZ3nI7R3NujpZgs6jcadT7UzaBN1ZLhGV2CRmRpJuAFrsk3rXh
tpRHC3eEjXdXqtkza0ib994pLQD6dNOrauGoKmRn6GdUS5TeKK1XLrQP6RD8dMkP
GZIZlwpzD6dLFXKGUaYeMYne9it+g457z4y39w/vN28xXl92MifQRrHC66FJzz+a
trc7TOvLuN4yrQD/UdZptywRDFz7ydi5eV9ZomeV8URYjJ3rCyIRfOpT3SlsaX9m
DQYsIDcDHjqWzbgHAdrt9/GOwI5bkpt2KviWB1/wckKzb+o2Cj8TGfEUy7Quqvte
cXwe1QMUAQSFXqHV6u00OU2SIPUBqj59FPXv+sHUSrkpMS0GyVMjNsadNCKThlRM
mdkUB1SeIXkejs+l8OqRdXDqbtVTN5H8xwLRb3I/z8ZaeDSprdhi2E+SYR18steC
wuqt1ZymqcTFoRVKYjGd5uaf9kFP6kLuEVjpPUykbHNV/dyiDhgf2Un8d+CpxREe
82Bx8I1JuvCMuXrhJxEr6YUV5YH4HDl6L/pn9fUlrggFsTdM95+WMjwq/hvM43JS
dmDnxBtQfI06sh4fw/GB9qcMtLTKVqF53ZiMm+rllu+e5wQj3k7bUdI/Cd3IWVoO
juHjja3ZQM5/KizhfknZqfECGqt+/UL+avq6ASAVwes2045K3GSh3ZgRvDj9vlfb
+rCfvseh0fpGVbOQ7J5mYsvF1n8MgpisBv0pMiAYY15Y4dQQ8EatedUK8fkyPAIm
87jADBz2aF5psNg4fwuhJ7JtewSiUR1GVxwjQi38I9a5M2mUJ6Bf0kkHNuKHCEqn
8+Oh0YeMS6KFKoEM3eTAOlFJuhW3L9nVeVyV4fbLJZNlwBwM9jLGIUNkTRB8Wkcc
m51fA4pb2650nMo1dj/CD+I+LG52CeaHaVwiA/dhKUhTAkvBi0b2GCFdrHeVhMQD
eERdVDZEd8TZamGPYTed0qV13VVoY2l5suBzLE/URk92cU48kndL//f4uLIgsBSL
smXbvAf6z+99/qLz+Ska2goG54rasJ4RQHxAIEvgdP1tNV9cuDPIfwmfu9Gqoid9
Ic5Mb70Gl1my60YxyQxPxJJyfrd4otkdXgdyo2sb0ZEY87TqExXA8NChnzHvI0FQ
cb7HyWZRNKwxuZp64w9yvlw1SiybHIGg0l7/nQCNFBfyW/9allw0AyLuwy2WHL48
GSi4OjlGtG+v6ApDF/UqahR3zFWUCmpxgwoMctXhJymDfaxhsLWEJXN6mTcShiji
EO5fc4BNpNkjx6X5RtCUJh4Tuqh0GyWP9BbQBdLvkOvgeceFveXfLDD93crWpdfb
AmZkZUNBbdxhpkdE8o9/hDb0VAZZrfj24GX7X93NWentBA8J0S8PL76vZ8NA8DkE
IyDS0wYaPcbpzGzQogcZmkRKw2s1cFENcaCkOjnXTYl/BmX4Dz34ZT8coKuBCB5d
Oxz09OCj+xwM2ULmKV32TXuY704IC0J8tR06PNUPB4THHncptOfWEETM7eDfPiVD
0kGPD5986dFTHmNPqelDJPrtgAsasAQ6Eof36bIao71tmOql4pV3EGPMEYQSWgub
7GJlSJRUYU2mjosVqPYUKLHWbnjyMcFh0/z+KIJG/5cYtWO5InwouaYgUBH+7mre
PGXPJmAr/+/Lbda6X99UAzTAzUDE60CUdGn41APeBZcs9i5qdfcPlwlSC6o2r0fD
VaynLs/gQJUCCNuA3fwvB7dkrw+ZyadI4zO3/68YQgSyl/cVy9JEwSi8BlLh0oaR
Z9FLKlGAi9yDwmd9zoWCiAswkRVRhfPrD55R/kRv5FgfaOxeYr2j6U2rxd2XnXod
y7eSdfdCSAUQjVRiRG+fTarBm9Gdme2jEwb6QOcWJp6eFtKuE2ekVfgAmauwRGnT
j9TU5BFwCEat3qICDrkZ0N00c0CucWSPEtz8CSy6rcoP1DY5mntSNVEFaWP+3nA9
VNH0aG4Z0lg2IScdzB8c5VrTQEtFYxanSvTMME9XkNCZPyU4Kyx/qq6HtIafxJz/
XIvVAo7JQ6VsrH76ffTOt0nfZpjET9S17nCCQ4pv7Uxg0Y64i+AYmDdkLjXba1wE
MBjWoftjnSeuNDraNYQ4ZesQUfZnz2TsF/S7FO+I3ibFoo3ZACQmxf+OikhwMYtw
bUHrETWJwk/H11QCzz6TkHNnhY9IKYQ/f0LUzXbgbFC5bYAUhILZk/CUnXsZJ641
qmPHqzo/FoQUrKFkQKtmHopRuMmtL+M2diZyLA3SSW+delqZrkJNdqamsKjj4V6C
XxNzd1wSseYVkwPs5EVmta3hTCdXkT4uFRa7pFJirKF0jpqUIuOEq14WlylPO7em
UM8p/yKq/hFd3fv4wpyLeMkc73yCzHgBvRFArjasSqrSKxosxEXOvY/5fv1zLFUu
Psw0MUDR7GLMgk19KzOn4nf5bwCLg/ka8Yp0OFNK9C/F4A+mGqfLx1035J73MFgf
tCLG1UJkCoV5rToidz0EFgxf74Q5l6rmUq3Oh3p6h+JwtbcpNYdRfuQmhagkX9LJ
jx4cO18LFBKT/L8p5Vp8VCDApE/eesRO/dyqG30QEW3oCPX+o+pzDKxSeiQsTwVs
zmcNizy75EouWBzcFmWt32S/Q4PVn4pnXig+J7tzfQ0ZbYKfHaqk7QQoy78epvYP
DLNUWowJnhHtUQeC71PI8IkzxelF3xMBEQTwYkqp+ZWdxh5CogAv4blRoJUGywwZ
JqgXJsPGvjZUGwzS+N/hbdr33LfzXHRB27QEsOZTWeDt4+oHxbIcWCRskrmQL182
OhyVg9cCRHmrQWx/goKpS9NT2ZBq+e/NbhghweEII2wqlwycdiIvtEKbzefDd57Y
0/s2OpjYgdEm01JP8gtYD9A/niQ65BJwDGdkALybmxeQOVhalZQ6+OnuU/HAsIDu
jj4A1QVOtcnD2bWV18dn+alnQUszUhJF8rMId2WP+yaL7Yr/EjAkwoi1i57X4oiD
aOAMAEONuzlDEEz7XALn5O1wr4IPiHz8OgHNe/MadSvcKfXxrWxPHVKu3DI9sxX1
hCBKyCuxRm/mPsLDZD8lTQSKJ6GObh4Q/FRdsf1pttW8AppXC9EiNFGtIK+Sp6Nu
LWE7MoZnmek9pzqp48/1cfJaBBhl+T2pC0v6KpW64ohh06xwePE9awp+iMy9Gdt9
/UIlMtwifvGftd9R9laVjqFOgd4YeRIm7AFAw8lwBaHQwoA73YP74VF4PdfklHAU
71zd+ecW/FlZNVYrk9F5aaOl2cRFa/zXiIpgFSM4tKJBS3mBObDrdDK7pwhi/a8W
T+8HZX6l5VmqGha9h7X2r3gXYjXXZ4tlQjweNtl7RwY2rjWC7TvkvXldt74Z18O4
Q6aneJu3hCyHGoDsL++w34OkUToxcwKunjAwwyiHt445tMAyrNAngGqrYNw+TyHL
eb0Vh19hNLGyaIUH4YDEtt9XVc7SnJYmHCuPRxSq3K0y5q19Ffyq/p9PS65UK0eS
s6wscDn3r1xMOPOsDuFzBxGpue0Q64h+CE+nAdlJ4U+YdCgDqchhjmIWvGZHQwRd
f8aZyS+k2zaF9rizkdjLVBjxVKaBeYMq830oupg2pDeq+zgfWXuJgwraxw2gbuDH
ZS017nlHL/TL2aSdCtY4bkt8yJnusbofgVSVi8vMiZVFrgDdWeojRWyAEtJtHhId
CdhPk8oONDw+UPrxwIm0P8Yud7iKPQU7GZ1cUbtxmPtERH1JXd6BurZbrCvyN4cT
zxouYVU3AeHoqofqWXN9etXWJfF7bLWuer+LYF3iDVaDeo14Xvg03YDPbfywKnkQ
9lEifOz7xNLZiBrCnxoem4nWbM+a9ALqG/INRuSiEMtxFdQap3F113WuJQdS4q0R
i3hpwS/a9l2IaZvoh6pchcupnsc4TxzfdXZaOEUj/tri1uZD/dWoxglM7ivloU2P
Nh7GT86K0M0n7dpHhdogRnVxy5HMiGaVAQTbAa0IpB5d4LItlouoRKIOhEooCJb+
GX+0gnB8Vg/LysQjPZp7unooNKPyNkj+3f6Nr87wVmdBuLntG9vFBHbad0YtNSg/
tO2cn2BTeTb/Yk+lXLVMS4Nl21g1MuExUdVkdxTuZ/V+36UqAYToNW4ba/Yr3I0n
VA1ghXz6czndEWqOA4k5KwjuTNZcPRKYEgq37ehVs7Znu/Y1OWNtO4nGgY3Iamet
AYqYtPLUX6Qb4kt891BRrrCPosze0KPHzuJzEEn5dAdZft5kdQQ4p1j005VvZXGm
85pqCPxGK2omSB1NBwhlHAs7SPjNYVef2RoP+vA/OE0DpJLSgnguRg0O9hsH6QbO
GgYlGDJyn6l95pM665TQ9OE53VvYAIC35MbfAwXPBB+Axm0er7H4wrWdqIY/Ar7W
8WuNnhTjtCYyPOJn2fN5zC6y44n0j5MhxK2bhZM2BbpqGvAJxrZMJPcPnM+KgTA9
Rh89k6AifKGC2i2nXSPAJQjjsDlqelkiJ4NNow+MtZt4kmZ1CZF6MDk4lI7qKBCS
IsbXTQoWTcXIWTYCJnfS/dCdhkmYXprZYFTWpxHkMB44uU0/FqgjsACDkBYyIm83
wNuFz+K1GD/GqPyA+vdSF6CnhAsG5Ag0Q7ueEoIQep3JYZr5A9zOMGs8QvqZni9q
TqKFq2LvVwljhvEUUUGLcUJ4AZIzFLjjIzrZwN2SGwkGsVEIN7O+IgzrzzUEcBJa
RCGuObaTxyYu+6R71aZ3W5x7rJIBSyywLZN+taL+QCG1M1z3yGup+ezGoxzQnWI3
aKU6cgs0o/XuUqgooG6hXtlaEJ5XLZ5LAa8ZdjxQ0MG220wPDXEbWzYm4rlYD88p
Kf8+9y7r0gxLaZz9eabenIYrZmhfCvwhZLrnpcotVhLvdAco0OKElRfcMjUPW7aH
UG64RLKk0AYQVpVYI7wcqkPAgVD7NDBy0IjfITLa7FSbrbgqLH5n3u3ph+/aU4vf
9XLia4LVxbj6ghc5iy6E3XyS+KHYBlc2Uz/jcyxTF3F1rqAqzoVPx0iKRkW08o0j
a15boeqbk2rQq7l6H51K75qzva3i/jRlIZxQ45eOUSlg/t1h9VjYKsX9sCrGwrKQ
PLIU6KZtSdiwnmYEQfCVfxKecSDvyVr4nXON7d1Jz4gBomo2aLr+DhK1ueqojjf/
hHKz6nWd8TcUeXTUOFeVQD4b7bd1L+wISjh22A1tFpRu68q2x23LNoZZw25BQL/d
0ClIf4+m3CK/9Fp6DDRBOqiCCV9ypdKR+BbKRAyTlFob/esejuzgaB0EvuwLRxxa
SQkIbUTvrWvVFvDWc/DwNAPB+hKtl77GwF2OgdichVhMdBIuYKj8E0KmxDknqPk5
5OxqZPZLSmC0URUK0bxYzYft8SvlBxzQDarhCiBZUoKSD+nVD2SHZ5N/iCOVcCss
V1P5NV8ldmpwKjxm4KJN4mYG3ttaVMOIgss4dgbky2o/Qb495puL574UBwp0yCsE
hiBT9XRQ7xmXVJf47ShMdjWb2Q29XeIDyCNvuVHtxje9N5HD/iLQ3qEYqD+1zc9A
GtijS/F5xzIvBZvWR1SYwKzhEkiEmgtbEu50XlD3S+XU3Tw7/j/nGDiJZi8n79G4
PrH/438eCraEa6Y10gybLPODuYwloprud7oJuwtTtGsGGlfXkgv1nP1Zk6GuxTw7
Ju6XOE3FVViImOaqLJChIKA324yWoeRe7CT6G0c4VRWnwO9Ol/a71d+eliJ5dkQ7
ztlZSyP9yAD/j3DvtysHdfDGeIUOov0mh5wXyuOUGwqMb62CmN+ml1e1XT6JbBbN
Z1Beh0+CgVEP163toXLh8fiJNi8M3GikMuUPSj+eRUSGjk2YKB0q01YTXFOdHKCQ
zNAfTjZtU+7CtHLVBCYXaFcopSj6ABFUvlmmANolKApo2q/xw3rGSQIPF3yJ+M7h
aTUqwIiH62vvCDnW3PzbIORm/AsZdh3vQTCGKBdeXwXQQLcLF3B9fXoi41ZV3F2O
wE/cMCEdB6JCql1YM9VdGj9fyxqyZWAbiycMXL9xNNvtAyInAg1068rbOJ15/prs
Z+ytzhRWJG8C+VGaAaxkSIWxpDqiEU6a0g9NFhgPluQUxC5RMgTkuI15O3V/49PY
sGcHGeNvRn912YotGy/+9kFMRMUDACIeMYxDsJ7zsvxDnuQxGk9v8Sa9f3W6/Igo
grtL1I+UUgu5aG4V4f3n3bgGhxZrFv1AWpgGnLIlVwS3gJxG/mZooITqFBd8vD56
BvWc+Sqf4b8YuzaZ88AHNrGG26JHBwOxvhhyBqEw8d4GU3gJoNRf4O645RCiXIKx
vgUuNruq7fqt2N9P1CHl2pkC4nDwzRWxXvUESM7x+4XC1dk0kS0KpPCwx4p1+0bN
zorY/S/Mphsu78+Xx/68/qKpdhPhHqPuaQpjjpwE1oDScJNr3ugExNBHZvScC934
q0fByADxnb012Pk0buXQheevm3F6w4rO6XVIyxd5RCs+A6+6+3LTJnaLGImCedri
5itgApFuvJ6AMdWWT4SekO89vLp1nhf3ygu2lNeSUQ84MDiEOd9Xpa69AKcN09uv
aHxchKu2hbJIzvAl0HfGy1fw/waS2jR6tzNpjV9Cn6HwkBgo19oUTS/USPmbnaiR
iBjLASSdstQMeZxu9JIC4ZbPXR0IefMJWqROPL2foQ2AxnyJ1Y/S3SUY/l6sT80B
HIU0RPNGm9didiSAdhhUly3jXJnwas8vDSs0ngdctiDllyntSOme1WTVomSu3QDy
3fOTsWkAcvTfhNhvA0WolfE9sP3vwkzpOUJjIgUotCQaSCqigPN8YSzsSwki2I+n
m3j3vmp0x4vNjdFBmq3GX7p76ByHVFS9igGB1rdAah/Q3TW+WqRCyFnx6jge1gC4
HBDcxoZmMK4V4b/j9Pe+T7dnkerbAfT9hmFLs9LK5Btx03HmYwo+Td3YrupNxWMB
Za+3SyYUj80YzqGCorL2U7taWUCQjMCP70gO+0/XIEs/PgzK17ygYeGn/RkN5Vji
7zVXdSTTlEWXQoqNJoAWm9VLLiVGCCzn9C6Fltp50ZvmA/PZncIzjxlTeXoIVAeQ
K7KdNWy5AHfmOoGzSL2bgf4C6eXYExNMxxuG96YBUmJNFJse+fyXRdTBG3mtY7Lq
DMZDCvOOT/q3pDfAXXiycNngx4aZwPXjVT0qgn90oYWwQsuK5WV4z3uDhu5te3SU
+HjNmnpLs/4weOKwr8K9ugP1SwLyNEQeZq9R+5iL+uIiPzzlc8yilhwzUYFpBIMG
RQHyUmdPrDWm1pRbill4mhSakegVIO2dRc7y5niIyBoZARaOWFnZu5ubBsdFTT6Y
emEIYp5zV0NM6IG4rDcvSPj9SSJYjSFGFTZb0epy5xe/t8Buwv97YHYNR6ChQY4q
4mQtMnJgux7r9cGW1LbASwuuYB9xqwQTeS4Z00QxEL07GiC1m36GUImf3njXpgYp
ks6KutW9y1MTP5fOGY32kQmy234k/d/nV593PDaJIV3KpSxoprAaiWMqh0GtTvBp
aedbGHZf6PI/hA0DgygI67yKSycVsMEfUAJZJ40KrZaKHvF/hxVNlMUc/P95qQW9
5tIEphmCjpjCCUBkKX/9rxdSBRShBp2lOKYKZhZEbS01Z6297C5AOBCyl9AnchlQ
eANa1HwSSBEieX6dL7DghWqShTj2+vzU05DYdXZBgvIaPGfk1xSDHt/WNIDuS2+Y
TDw4rFSjFiYbAZOuW6MLTSsVOwgYwoViZCdesxKqNT5YMpKA4psuCx/EMLS0G8W1
qc0A89+S5IISJjOZj3TwNmRnj72aCYshGzEYzwzxxqHPdkeQOFNXaqulZztaDsX5
W7X9lKM0p+jqbJiKorbCDPaDlDDYYKmepCwdC1jCCTP2yn84xUIZvpWUZYrTQNz3
n9TfISTPZcxT0rm9mU4P9+5kBaW3Syw3l7K5VOhT/zidlKnHbo4e6A4G46ReqP22
9/xw1J/IYJDfwxTicOOkyLX+iM1VYdEbeNAnPN0598qbiNHf55ihs0ARlRkO1ei3
gFSWYLudVuVAF7CaeD32t//94FqqR4M1czvBw7mGJP+ypHaE9PxFQDh2nVkoOVR/
k96bEmGhTY8LLPp1hDmt1lDClIx4SvArjvluV1STi5UGZH6KI7ZBnbFvYZ7q36ss
zUsKe7A0Fx46giy7Z0WGqN/inLJSyUeGMM4/ttyiJVMfaWRJFiKqCKieBMxKnKy9
iSRMcp91sEBhAK8g6Hh4Tojp1hlomhnc2DtMjkQNl14HqPXhT74Ziikkl6p24Sih
U7O4eHXwrmwoGHy3n3S8KUd2f8OzeWaIJ8sQYsXozvAJeMJ4SsWpN5n53vXukmf7
aG9LEjQQJW6H/i8VwQ/+cvgFCGNvYzcAL1sRn9azxxRTo+veexjP5Kge/19qxQJH
AJ7Ie9pIKve2fA144jq98nfyYnW0punMFzQ5PH/FI8npsu99ksrcQqDtG2RXCfWt
UAVkjSftL8A7lS32igbFjzF7mdvjVORgED3ey2SEcU4HZYQPhs8tKoBiANc9kC/r
kxZQ3vrlIfUFX6yNAYMEEA7NUOti0DfwGut2xulaBEY+jBETnDalo9NVYrec3Ytb
1Re9i9dNGzmTB7ox4V31h6WSudl80Q9nJH0GCAlzU5Jaw1l/sXPlHcMmF0J+GU+B
afICXIakJDcjfhy8JF/JDsTlj9344YwFIrfDS7OCHuu/5CFblik6v+rOaEMaVRoS
M+eUbjywo7emmT9SCEAEN14YLlB8M6nqrJK/aWEyJua24Fct7G5aY5hxSyOJZ/Ys
gcJJYI5AVbML6mtwmPce/LtxxOWljt3sAQyXequM48FurRPZ8loN3qye1prAg6Bg
oXQouWgZxoEC0G+runhdcvGOLZO0zC063lUVtF5AYQGkt0gqUBh5rv3CFSYNNdxF
5gk5JnCeV7JGWyzllOqPHbRuOHVFib8Bk/aaKYW27Xcrx5IgqPCcf5DDSNCnpr5u
xu71InMGWvwZoqKIh27PrV1CUwJepLCds/Uh7Vwht6G0b/w9ZalVapUCPHbdK+1W
AYA2tGADuWzp/eDe/hB/d3/SJihfbmASikSt8o78HxgQcYvs1PZnfFQ+XFjYOgzz
c2sCCXWIlRcTUkmbqsHDFmhJ6jBv5Of68BnwHdVwkmNuvjj+Ka2kCRDNK/29wtZn
8Ly5d967WamqqgGz5TacKCJnlYhCFvTdlxweirdA3+D341+e/ADsi1POwyQAXdFX
Hi5sNBXH9OMaX9f3BcsWk0w/QwvaqrsJKa9s9LC3kaN6I8DEZBPpS19Qtq6hWBH2
3VmT4B2jTSTc8ALHkN8sM2jvvvE3rSjyMzHOzLEEgxsUUb2bF7mJpLbjnbc9Swxc
VRQO9aWfyldkdqK+enmvTxUlGIWMoO/xs8TnjDzubzdh4TMjytXLLqKXsSGGbAxN
UiM6ZARg8+BILsGiGxwCX7AVjLRuu4rAEcBHgMOqN9Xnf6h5a3m3iii1IKlQutne
1pqbn9u/Kr0FkcEkdk4q31oXsy9Sk8VGOtSctu2pTc26CtH8S0qB2wMlRSbCGK3e
UPCE4G+4sfJR5odxFrQwOOnOIi7kFEicVRQRu6PdFIPlR19pPf6wJgr/BTkjQUAQ
1j8q8dC53rlBMn3qxUTaNzrqMgZK26G5SCYbqt02mSLn04fRLudUZNWz75gHD1i/
wsMEybcZh06OAWIMioXxNAz0a1J87zEQJT0Ot7DeC2bMnhAnA2N0KYdsab/q/xyT
Fawo8LPZNfE9jbWhZXbx5YcNG3FKV0iGBR65Gcjeqj8LfHJCqtt7y7V/MDv5XqKe
vex1KP+FQg7mUZLJS1Xx5Fl8Z1VN83SSOff4fsmcppChHityVfhwJ9hmdW4fX4rT
vWrAOV8PWY1EZOAJGWIMk+C4T4pQt3/jsKbQpd+MVs3Ds9ypLfENun8ThiKI+Gbj
SIl71FJQPv4hJT/2vyA2E/qwM/NfZ74qEtPBKjfHX2iwDRJjsPIQ5JxsK06lFPz0
BMmB1wX2fbn/2eKHrwnOSPdx/CI50PqU1woGFe2Jc6AnKpBZyDnUAJ53IhsxEuW8
xJjlRXBc5MoZuMXKFCDlTbF15vxbccgOo8w+appEj0ARzNt8+kiz9/9NKft/ufnh
IKT6vuBSC3qYB5smUEYYuby0TJDUZbdm0vx94Kp3qRaRdhDwD27HkodH65mWGug/
BmHWqDTAIPrLB3pPduwDUmOY/BIEiKEJ6wk8OckjDkkQcZajL8N2CRLTvuPUX6Uz
ImkvpDaoTd90/UxpcVYgeNj6zlPqVyQm67v6gMGiTscHcFDDovJzmLnyoBLurcgf
k5bq2T0eMgagVwKT4jDKLej1ofw/LYJ4zw9clNIpWDtNa1P5kSmkqyCO50wgfj+x
YnINjwazLNYAb7yoBagPTIGImLKBNYBJcTOeiHR+XzbNputO0XpFEt0EAKWdCnQl
r41D0Xh+jmDRquoNA36JrtKp6OeQBJY6Y7nMSljFF06bHEhHCrYuXj7swgVjN89d
MMn9xnGFSl7yI7XIx59O8Jp5OSSZMRj+8543qCnlGzgHqOBmFKNR5dsoSHEZ4G0P
/2QQvtTgL91iPQL7F2XVsDCo6VXaBaiywDfyFosQcpP2riB59yoa5XyJPklpserd
4/NcVV0CJbiHS2RxF2y11Kuh27pi1UonWZnYejjTny8+lCP9tl9nMexoq+QcjLs9
IKq4xk17FQQFr06uTpxnZEvNFUTZfFViP3drVNfGJarbKm8tNcp0vqVwkgRvnQ4H
qq76uz5Bd4F0i11cfyuKFoha/qWM7VamWmlpju8le3kgPQMSgQ0/H/TdheAQs2wb
TXU3P2b8z9ZzPc7OjUchO7CFJwLbmChaWngED9yf4gmGyJdpRPClmB76zhWgcE7C
9VYjaGVVNULOoygawaOrbGR3SeSMCBV+cXRaRh2lXbkMLuDcQHGscLWnQwmiEkOU
CuVG34wi1B9reM9OT4nl5alIpS69xa3Eqix+sG0qY1VtpfGIMCFKZU29IqN1kgY4
Ayx8cjBw1zjPhMyuYHUSct87VM+aPDfhx3RZCPU+6A8nhgG3DsuYaiHRhvoZAkEC
3OsZKlsGfNCB96p9QM+cANQlOfHW4wbZAdvwLFP3/w2EbgWC2Gjjmdk7Nw/DkNoB
G6akGSEVlPeozwdWBzHkqy1tSs7GO6NixH8F+C10JrtUEw+cAXWsCKmNIWd1vs8t
pmO4IpBkm29HbCmsupmcmwiFijmQH9EFc3EaF5FzI2r486b/lHwj9vACqbkPU9Wn
sXJzf2IHy9z/Yh6CRO/YzFD1XyKAAFPoVkxPvYesyj+xSSpRrJGqGg2CetKF1lLE
hocokDDPc1JZbUKlR4WRJz/49ZPUWyFYTc1RDOEVY/Qk64ZS9/KHKlCGYuz+n/iO
jWFjH5dcT8UG76Y5ibh9A77hlnxyXo9PEc+42a/QVwBdrDkzF52zNlsKB5/Voh5Z
0zSGgSWe3LSkaYvDMdQnuVlQiUld/vWdwG4qKPIfy+vPl+6xGnreMicsPbkqnJ1F
+TwIXe6fDaiheMjeXC0X2rV4PfPnnIhg8az/7Zrq6cvbmE+KFCj3wfO6kXome4oy
V/MXtPkcJ3yVZWXZxOduNnk2ztGUl6d4djKxoiVGUR4Edj+ujCo0CeQauSyfoRXt
jR//LhEHslH+ntw7AalfDSAXB5E9lLmZK96LVehBRgjBAzfKA8+6IN7rdC9RPnv3
SC9wz17c2EGIooKWHrrzCw39A9C2dP2DxqGH1R9ZAx+atjafDHaR6JJ2U1/hGhYf
+XBjArqBCzfeZfZ66WG7ubii/ZQkOzTalfoNCi6HlE8/F3LG4ifw+GBTZmmWli0e
3oBJiHZP9eKy5++vbz056OZTgK81YYp4PJLGMY+k219NAQxVzv7TUuRQt4+ZP96K
SfFJxcrEI8nPmAiSYErsLGxfW8B0LQ+Gz3gTDL9ujnp4NmYP1foLS05udwfiLWaJ
SeJTYd7lndQ8I5viuFLeS6vGSiPeZuL4cMqaYDcINMbjrMLxsh2tNZSgqUPCc/gm
0buSKbi1KgPBUUyiJBugBx/1eofwBaRHkIs0UwrY4pvuWCyGQXpGhZknw7NTWPms
iyMwX6cvGfvUdYBeKuFO9Mmbj+JkpDH2FjE+aLUH9oO4i/5XYEhGEmQ9h7VxV/rs
D3tQA+VZ/jdq4TErSqbFQ4yHW1fqVdpmqJtI/RXJgFOsxxqyInDg8lN6z90L2gcM
8WcLkR/6E8j0ZV5dqNqhfl4WrDncCNWhpxP8cPV3EJ1nJB4VJcy1BU2qiu/IH8f8
eZ/xmIL+GmKlADZKQxlRxZHeKhILd/qLHETKQQKQBBU6mlWwa7f3nTLCnT22Hd62
1UpIqwMQbQ5nZ+iLcoB8/nG1+AV4eSMVyDqzhAmTS8CqIJ3dic4u5dkYQcq3fDkN
qkBCm54y1DDfXcpu913WaND6hwgklP1kcK4nM06suH5zJekivfP/DJ6X+DIAJ9vw
0WyTaTD7w3iSv+JAM12oyqJpkPhyQIUDjkABm699sQ84c68RLeZiR/cfqayxQcY1
+XFRDrhVTTe0RqxkZqEWNvjWWxjj6FnTjM2PqSg9LSOqkx8MzWok/OAdbY8+fVUl
yWzuqUzclgmrws82UaYQ5AsFh4QMy57BAEkUMHtWdMlTCcx7ZFaTc3dAdxf+qeEs
Wfco2Oq1ivCXtK5H7dI9kj5K4aZ09moZ+ecrm6dIzVAmuovzrU/UkMr5CLp46sxc
okgDukkyWCf4JXvviL5kk4QQqMfTybji/f1mDwjRSENYYz8CWX+LNQO+qgMf0Z1r
rlYOOzqkOt0gJCmYLkh0i8pZ4x1SBGLVW4Ddl6WEn1RyKtDnMUIFTswNERBFqbyr
ZwI507ZzrPJ9EEBrsabFan/F9AM3po2rB2AAZZ2NF5DVBnoz0NRBCjIjhP80OowT
S5tIVf7ZwiEOb90qLZKYwnTr4ib1dO4Scv5Xz35/aG+WyeWBOZEugMsu8sX2Z6RU
8k5PRaiX9tmYFPELP4SHZotFI9lB11vPsICAiYqAwanaMS0Qd61ZoPyBLIz9r3Ee
exxuTb5zuJCmKKmoqs3gF/DYhnbLmO7dblGSfiC4a0pYGbmvUlfMDzQpMQm8P7pA
oBZr/SoZSQ7+UpDZZrhDa9qKpLYCkopEc067L0yguxYuhYOSph33N+P/BMkx+gMQ
N2+ZRoBo+Pq5r2RiH6mVaJZQjq57EgQtAgTujFUHa8nz8MQisI9m1PhmVQUVoP41
orTZ8SfxpLHRHOGYDJ6oH/yVZ/c8d6NJ5stqf1/bKhXXELx4e3kdXk1fOOnaYflO
wvHDLfQUaZeUvysAfG2FXHt0C5SpEvB2Je/6A15K7fPnUKX6dSnBQ/hKJmRvu+qa
+DBK5di8pOvuBp5ElqK0gWM578BsOpMwmEZKT3sydYbzyIsdqu6DzIXCFpxR/ptk
tuboO7+J1GFPVwNTUqWs0w/pW4JPKTbxEHmO3nUb1e2eR+5MUrnsUSCcgMxWUDXu
GSEwcxi84Z5FzKKTRbaRFIVqr1PfkQ94kZY/GAWmvte5J9JhrE/w+QXIcU4Qjm6f
SYnxYFQqkLsNIBLKK8Q4mKbMtEqEMc15RQURBAwKFLQhgACq8iA4sgnu1y70O25H
NLmPN2YjccO4PYFd5Wuoqcdzx4yGxAuuq7n+pARfjWNE2cBdwN3h/w94bB3WoTSl
+2ByCXDvw7qmgPaBoLYV9R4/4FiOAjhKfclV3OWFjholY8WNDf74Q+Yln0+urB4N
S+T0WRFUE9fxtH277zomFXJ/Hp8BF6n+lUQy6jLtnwdVbYF8xYR7MxRmd+U4Xme6
SH/qkXNv4zlCX/STK14IuL42MbmnlpKVbI0+Azs2BfC/QsoZab1xeApqBMzXD7pn
nL++2JosI5+IfnByu6x/6Fahw6T8ajdG8/lWS44FvuA35UVM/6D/6TfNrDV6uoAx
edO1kqyINBsCHg4neC0zPc17oRSZGZBkkp3VtlYVlBYE7Ia9C256MEH0S6bWwdZK
hHec4G3rWhMEV96j4coFqxJg5CMjvFiFbUPEP8I1iLZwb//QCZdCMxMTgOKAK4qs
FyN+PfIp0fLrI8AUUjPO/pYBS4QicH9gD7JeQPWKIESqtiD2J6k4HmpHUhOqFTBv
RS0nOdgXnv0La8JYjkP6iksajrE/0uuoGuotzT66QcRvObUigkQ0xh7T0qkPH86y
VDFU5IWIvTWhIA30eGedFvMcXTr9/+ruPdKxanKolzuLSEpx3liCk3UfgtG3UZpK
1frQe3DL9u5IIPvjUPqBjklaabC+J579clLa4nxcX/5/ECxD5w9uASTsTSl//ZIx
7bBDzaYT+glhSyHiz7cmP2C1DN/QyXED4ULyi6cjKf6rPe2IvdzD8AOIxtpqVqZy
FM71D6CzBqFBRXo0Il0VD2lGaHoMQ4UQ1xAUnBG5UQHpN+wrtELA50YqWEsT8tHy
sj2MahetGwKa61kJiYGfJUKVUJ4BcB5We1LBzolScWhIJCM1B+Yn2NuK6Z6TbCe/
E4wy3901hWa1FeBjNnfie1NusjWM3QIt9Fu7zEtMVG+BpeI1zmEvhtCcMtr2ouCi
REwWP1lJvqqZEfR8Q79GPOUWBVs9n97GXPg12l0HP4X5GciYep295Mnrd77mhrtx
hkJx64vbVPYiGutZQAFbRoh0GUi9+5KJ5q6oSVIvqN4Vev/Rsi2yyeHSUD3Z0FhV
d1ubjKtKEuCprlTasZPVe5dVqOTdgnMK2Lsb//15bMci6YRqO1m5Z6NLzmN28qlY
BbIpNco7NuJs3CwEW0e4xye8qEyx8Fcmx4hEBsYHpmzAPLxJR18ly/oo4F5m0Gj0
43fn+dhDlagc73NmfoKrhXpUPp4filkYlfJnIbywmcYTPR1nJN4l8en9O9ojQ2VG
wWbuiDAhsc51CXxRzDo0DTB4T1zA9dfbaRasc8NCL+hzttCMOefJK5INibJw8R2z
5Xa0BtCvyLLR59NPhD7c8F/ocjU3kO110JMeQftozHt/yxXSdfapQ6z904dC+6Zi
LibZytD12cEuMWkfqVnHugPzwAuWbjtdJA0lhELrP0rtjyC9KuKzKZarTYZTz9au
dXkeWso4M2D8laQHweevpVmdA5k9IspoTTw9cIjTewg94qXVXc9DRv7KuyRmxkC9
SskwbEMGS4zkLCMHBRIuINgRJc0ApnaQe7Z4tQ6ICIHGEURk389yRAT+eks58xyw
rp/ErN5yFP8Epz4uN/OzXxbR4RnPz2mludssVDa0GjFljSoU492Sg1AF63sNporq
rkO/0jCSgIq91XMeh2NFPrPI447UiveiLD/AdFWBMGl+uSEC8Vs+K0Zu/LI/5Ec1
lKJByFKM83/kJNg74e3Yk3Ysbtd8rJPZ1itpGmir1r4wWh9ZHnSnPxpIl70ZVDiy
YKjpoQ4wGQdaes6Q3f614bK+H42iipF8NXdXagJWqyVbYWSpukDoWt6m7h4PMh7O
RT/W5REGEnhgsaunm8+W/+N3O47167/cbIhmsTi2sXJ+TBNXiqkuSXxAetse5S+D
RiI2Xm9J6YSI4L6ZPyG0cXYzK8/TgnvgtsLDFMeSFDcQkAejkrOMIf3cB4lYs6mD
mRloGI1JwreTO3/Q5evTcs0WGz2e2a/IcOiHSNIpQDCkXvDRR8ftyXcgug4utayn
XEfJsIB86RQLIrht2qcgVz86ywD2d0YUMzQYQHAQok7mJlzUDe5O4jkIuRx2xcJU
zKMozMKf5Uu1CKnJ/AZ9RnCjukrSqZOmrycr0psNYKsPohUTlu1f+SKIheVRqCm5
bd3KpFMw58JYFZtKFDxpShrZbuAQkq/A8w5Hwd33g+NycKJUFdm8m8TX9eUKSjRd
eom+LDK9HIBeA6KRh6gJIn6K8nf9vByXxxrTCwhMGE3zlRLFoY8s1YsF9jY3RLxh
Rw253xHDPYO3fP9/Gjr1X/J66+l2wvE19oAa05cFKx0LUZpMWrhYKTJl/kWktYW9
FGQpe8AVWtBWFN/mTs4St4MnNaAoJbx/sOc6W/qiKDmyzTJc8eL3FKwE5VJg38Uv
iOcIQMJc1PX+kFj48TaWjKCEiKm0BDlWop32IKttV+nDcIw24XdnItiAfRszDHF5
zOt3cDOYlZOorl//QVCOQ7LsUDYYApjTZtTbLJrMFiZO37hhhrP2ommCmeH7lP9Y
ZaUJcpDFap6HCje61oxKwY5Xthxgmt8WcOLb+0/s+5hPdDlw/0B89A7VUzmMBrI+
EVxvS/c+OXGco94li/RrT2PLg0E0csK7pLHTITCN5y6FP4EwpxdmCTo8CbjpAQZa
aeMbABbQTQvIEpS3jQXdV6lkRaGl45h2upzoSsdvSO32womQVVC770dA+HAMEZGJ
2XiGdo2Pgd7SAU3XHMee4IScnirXBPIo+ZSCuP8QrOPuHLPmM7zgJhktE7c0Je+Y
ya/fVQ8sQ2dX/moTF+AkvWOFIENCIKAr6C/qpVZJmQdQI47f9TZf53vIqczB0jA8
H4Rz/OimSdFiYHzF5EZ0Wpr3umONNKm/nUwJKH8pQ3Yj/B0EZr64F0hAcAGf3j6z
saKzbspogPh2E9MTwr/DS0FbYoYCEQPD5ymO6mJnSbdtb1XA7/2cL5JwiFQ7qg+9
EjDZ28fpV2WUkwgLg65QM68PN5ygq5YyYr6nxZMtQ+cEnElqlMmjJQ7Kb3yeKUzx
eIk8jpIuKnOx5y3jJnIgoqHcbtuLPM1ZFwcq5xSIOxoPO1Ask8Ym4Zf6+OXLWFL4
c46G1VCRmgTb8XTIfY7wvztHl0Wngqih03h9fXGOreeDPXikz4ZChT+dQj6iITkX
3MVtL749pVzlblZSRtlcCH4NcJ5xgTaOv1TX2uwSY03uIwOQL3ECin+vg9+54KNm
2lhllTm3tiA05jigQ/ric7oWCxVnVJcM1BStVQ2UGM+U4EHmsSz2SrdSZxQnsL30
erUp/M9NyFY+Mu5zXM0gL1fQjpC2pIHPQPY9TUZNvEZ9wzBXXd6sell4+eYn6NwL
2VD1fZQzHJRkvxapJyucldbo3hpwxLj9i+MHMuXxHTB8Tk3674xoEn+g6BGR83+t
TI/le1pZFqOIN1nljt5A8Q/cohSCOYZUZgvIbuId94aEYxU51bJAYOuxMcjeyNAN
/V28ewOQmxErng5hfYmZcmGAUhKZW7IZveXmIirm0xQRpowWbbZsThcychfpLDu6
l/wWZo/LcX99duue9g8uBUe9dxzF1TNNChpZhWGj9m5JFo8p34nwb0dttd64Jdh9
35sBvL0BD18vC3XJDUICcaEhPT4jPyj7usJGcc5LUXnYwzA+HBce6iuhcaTHksjZ
QWSEBrfoAob2WpoyaKVAwtBw8xzd5siXVzrhBT4BPzKiiztPK8D9P+A1R3vrwaXt
oSi+r+ZRFmxbnZmDE4njLLnXecj20JIZ870WZTUuimiawLTLOfqC6dMmiuB+jHEj
2AxYGoG+d06j85eFnsx4dXDmrUw9RzH2EFfQqdxJ7iH5+6vtbSA2kPXSED9o1jkJ
3HXp0Way2gjCs7YhmZbSrMWlmjjxIvnCPPO5vQlXOiD9BLdQN3Mhga8Tmpdcb7tN
I7lxkUOww0ewfnb6bKR/6aDrhy6nrEt19HMEnYpMBsh8BC3+hV4MF8B2Wiq9bu2q
PPgQ2Et0maClFxmSy6hg0IBDZb2MrJNpOJ/Kyb5STMkykL7jTwqfw7qazxAsg7TY
U8X6ivBj8xMdK2Bz+ssY/6rwxU4OBCVWADliXrASKFLcd1ocFcx12h8jtH0e2KwB
ftEqoi8bI+dgcwW1lLdBBWIlhe/z3bcuTt1nqfXyONTkny1n4Z9gHf0yYreg2moE
ncHLd1LsfS66UCYWFZ+adn6CMXyDH+jTVgS1i3BsqJGrXueZdzteGa3z1GIRsx+m
oLYAq2JIxfNsY4X5M7IEOryaVQhmK5+9TX5C/EIEZHjfCMAlvC02kLpas7x8jrUe
8zt8ZrwvRSS33oH5lF75NKeqYgkoDbJUFe0yi1dq2aIJUBjK9VGW3q3Hg2qRvXZV
kCCLJmyqvftcrDUA9iCi866ZEiiDirgtBfaATN52GJ6nwWMeOHYmmK108xEIp9kY
O937JyxqtwV2dAqIkFtprSbF4i3oqai20Dv+knPpLRzyP/8RxxOroqWukEACIldc
RXK1nW4Cp2NK3HVvDRT5R9Do3Hk83ojAKO8QCIoeb3XKSQkEJirQGvFgDd5II3v4
I6JHCpWeNdOouLgFKqfy/KybmTjPsTNVf8UvmIBbFJJbswuUueUHQT8iIMoxrUKk
TXNRoXoIxYMGK/+Ph78715ySb4AF2MnKRm+ufC+poVNNUuz8HqxodNjK8SQ8hLxW
4dbKuj0HD1+99ZmM242mrSlNMsgbTdRZRvcNFY8BdRyVpKyyRr1CznY+S5T+Zy+R
ll0Urxzy9VLLl7Y5cNXmNJImA0NsuZwZeahztYZRbdD/b0m7pDsXxurHJHgofaGp
fCGxv/Wml1hnORhGc3wg+OWG8d27ZdhuyVbMSAe9pKWoG4UQyUl9ScfGwkPSqVWW
Kmyr8v2glfXk00KIEhe2lkPrERP80fYDefw6Z5IH6YChaFg5lTkppGjI2uYd79e0
ABKuaXB16GJU/8lSO3LyyrcRLhjOsPIQ+S3tA1xWFg6/QLglzzwHfVTc4jq+01vG
JJHqFdm94+DrUIidsRlMfaJ66L1cDKtEH1gmmxc+I8ZQ9oHLp0KYSEAJLIC3aeNg
PLc2RFR2vpjLaZYUZRQA4AxcE5bXmdtItwDxyw6aUyZ/mFD8a0oI8TpSvsAojhKb
BcLSRqVGEHaRBfvuiPkXYSASfLemziV47GJC1V1qnjkw0OkOwvc96cOl60q7/X3r
OlHYjNnK+5TUTC1LeYlZCpQmOFXqmIOJpRrlzzBs9cZjCfXgsl61CWOY6QxxgKSm
OrzFtLsDMEyRZHZhoHAjUmvWFRAlipLsoWcH4BwAd9rP5fN5P/OmV+/xogHy7QaB
y7cCTstl72Kh/+R24nIoT3mfsfDsPyowawXdD7Isqe+yGJ7Jxw6ck++MH2rrGo85
Mlkreiz/czMS8wFSprDj1ZecRvNDuYpEk1OfAmDbptt+hf1P8Oh44xIMS9QKI2gt
BB3K4DEq1cDFKrcURmzHVGJ1m/vu2/s/T9kIwd7ZviGKCiZilqTyIjgFROE2fsp2
XWP2ekeke/t2kLk5YajFF2ffNgn5Ro8VBj28nSC5zPHUZ3DnDHSd2Xd6ac+lEfq0
CELqA6vtdWNEuSZk9NbEtKi+rM0nSBjFslOI5Vymv+dK6fXx7vkHSddf8dQNGSGx
zewHjAQnpApkvmWaQjbFqqyTW8FOkeZKtGK7jMNdcNcJp9G1HXziXSRWNSckjrcm
iionvOLfwtVHa1w+pqwbqkR0Q7PLp0r3a6GPMil+WmBOBese1PM4s6GdfyAXsgsY
QfnYkP1NQksYG7UMI/XECApO8xhfcO00csa5ZGIM2XY2x1gfPIkp4SiG2IErAIRM
sZM1lfQBadxZ5HdI+8C3vuA9VoGCGBmyNqmWqbnl8sPUujE5A4A61Pjflu6uJsYH
Kd16T3jYrdHpoEsqIfomqkooC3zWsLpd+0cryCSrDeEJxGwfD6qEEUS5+tjXAY+x
hl2LH0nzhdInHaw/T14RVNBp0/W1f6Ve8Hq9OCrmvbdhrEPNC8ile2DCgpPxljCG
6RX1ZRj6weB2I1unnmun0C2ER1Hat9ngnEUzOdUr8uA3XWB0B2WdiEPgP5y5o+Cp
NZqC/YAo1Gh725ZuMCEMBkjjNz6yq/3uqnJ6ReC4KMjbLnHUgSSpEykgH/qbIjQG
//pragma protect end_data_block
//pragma protect digest_block
cLZIylPeFY5utsLDZiwIWtJyDWU=
//pragma protect end_digest_block
//pragma protect end_protected
