module QUEEN(
    //Input Port
    clk,
    rst_n,

    in_valid,
    col,
    row,

    in_valid_num,
    in_num,

    out_valid,
    out,

    );

input               clk, rst_n, in_valid,in_valid_num;
input       [3:0]   col,row;
input       [2:0]   in_num;

output reg          out_valid;
output reg  [3:0]   out;

//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
c/2Ff1/3JO9SYMGXwUFpe/GVQc13YG1y+czvrwEcUZL/orQdZIam2pmIqxkhC4iM
8/UTKD8tUiAGFDfonKijavy20oPMls9scu2RYSexnYLVMZtuieHfz3NdyyQLkf82
zdjG7CzAowa2m5yuERFHQgUBfZLqFOn361TDG9VcJGbDHD5V9F55EsCZI8rRtPn2
qJWi2KO64JYlvIsvlKKcHkVucX4+C3vfpgHFZQePgd3xj/OhXr/+1mVs6gyGn7V1
rUQWs3ksZXtu37jhxA4ZT66OD32jCsYhlGHUVJ0aAaTE0WDWWE7spTWT/61715yA
gcHNx6CEFTrMMt7u0abCTA==
//pragma protect end_key_block
//pragma protect digest_block
2n5/AqK+c8prpEPi+5UeZ+L8knI=
//pragma protect end_digest_block
//pragma protect data_block
BFTzdlLezpjtykVTfUR/KSeZxIxHLLQViNLIg2MGQgu4LPm+TzziPYivi4taMNSa
vGntPjWTSaE4G4Y+vLCuJGMTvVzm6AeshK6OjiDlvpFaNFwW+w+tMFCuJSwpH4Mf
roD9g+XJjD2ytQcyVk57Z5fxCzYP+L5S1NM64sqZgFBsrA7lNUAGeGZXM4e2U4vZ
/q2S4RG9hdFgzas3IjuuCuK0l81IlOi8MRctD3Lc1pm9Qrb2dih2XUQAkE0aA8tX
RrgpxlI0BdGZqwipsdI2GDmxMJzdicHvu6IRlmSlU68FXZxmLIfbXkS9NNZNanhs
ZnFXmnxW9RUBC0udn/U12Veb2eMw3Idp6S3xk4A60lh4tB2F/0CyTu0hkMnq9Y1w
UFJ0L6lvhnoboz8HRdqzNhz6fI6VzIPTOwsOxo3ToHdF789MXSrZpeITqizRAZ7a
OTeUrhv6kq3i7LKUfL1s+ke91lBDPdoisfryIELoq1eYUOHN4k5Qm7PbOq8bJSYZ
mDN3VQyOBhgnPE4khQItSx5FIe3ltj6cXDJRSPDof6RKdtMtwH4hegwBVSqG68QP
V2en9KC9wjiaOX+ztizkMBGyfJZm3ctMs1RZZR1ImkNFwcTvHXoIt8MyzmzLq2sy
ZHsqtXUstEvPhbflw8cTgH2UrhR+L29qIWtg8prIb2UfcQzTan1H6dzaPSp9T5NA
PHZMfhFuPFTRrRGjNx+1b/fw3y6krReHsCfFg7GKATlXP/henV8oeTO6wROg+OLZ
9saaQ+E6C4JSvGQ7zzglmrV7zyZO21MaPpQigXXAXVwUl9XP1f1FGjCMkcqiErzp
Cd0pXTvfRDOu6L8dD4Vrm97qRQJ7XH4uKXDh12a+lCz3jxo3kS2LbLiIfqirkuwb
3uGfy5ZdBOlI4tT5op1HCWZMQf/OPzHd8CmMvfdLAM1OzZL9dXIeIZqsumpaE+Lp
t8SWtWiaa7MP9X4EBrftxCz6k5v4hvZ9o2tfY+lrTQ7r9aM5qLO5bpC494ahgjvg
08eYdIbwPnRNTZENsvNtPGiNKJ0Rg3PMtHG9VgfveUQTZBO4IeBoCgnyoi7N6/EB
HTtnWtAWrNSIlTzQWRi65X54soIwrUSWDtNbOV6XxS5DbKEx335WZwJkgwtkuUav
Ar/APAKKFThFGjFFjzFmOoSKKZXLhYdnj5m4hkN2Ozwg6KZdgXd9SXXOCGJTT/X2
0ZKOJIia48Yd2qkcPIapreXkgiT9y/S6/DHWTlMKpg9ouOBos3O6Dp/JUZwo98ZD
fWpF/nDamaip8uwW69QABodlao0uRxPqiL/z/IqNQ1hxKwWdRD6ZFUByKd/4rV+y
NExS72zThpt6/LXv75e5BQOtOd4zT0aO5lHeUjKYiEyEcFDVkUrnuyGi2a/+/tey
e+WK3RVR32mrV9ye/ebX/tzeXZZnUINbFrcH9sl5hwdfGal0wI0OuZYszuMqm/8w
BkANzYIyAqW0gXPJF2mXvR4BdpJrR8w0MoCrBbrmDsYUPCMV47fTLV4QaOGVzLKK
iz956cK8B7ezKCriXTdubwUFpWcE/D0+7HfRydrN+MIZYcS1RoQQXw3exNbwKURp
i8jk7wzogI1lfzArs5eGi+HzZqD5hpBvKaLb8QtPHWjjP0kitmYeuIMWp7vfCne8
Tsa3Zj7ueewmoYCIUIYbMavRAnFERimPbWxPQpzEAFuOK24SlLza8X2BIk4N7+Lz
0BNUvHG1H9v9WF+62D+p8PKc5Jsa3axaQpT2HgvX9/0NyFXxagJMPPJ6jgYab+Vj
g8z4VigT6Qrb8AzrPzOv9s5/DijRIg7mgGq6OehS3ygFvV8SZ66a5i43jDgHlFlS
wz+h2lMKzEb4sZGNEzynMboSfM+vXag0foTKifIkHiPOA/uwPQBHbPxtNqoO9wTk
jZ77xiWu7/q2m4SR6Mi1fCw8k7SYhpxizHCfXL5JWm84RDTaKWcbvgUtLQ20jDpG
S3lyZaEd4RG+Ok1gSAsPcVCqg0wKm1nk+x479iOKG0pkl8+u49/V25bd4XoJ5J+6
19si7ykdxQ4cFSPI1cIh5YXMDbUg4O+oMuOU8X90PfDfH/LwqDRi113v8TCAsnLL
BjMhetk5J69Q6UVP3u84qEjQ0Aln70rnjbMoqGoPvH+smipc8WfRcfoWz/+0Y3S5
Th6WXuMNOSaiFxSvN+REHmJ5U95MQNdyHLCh/SmhFsz4lXyr5zV07EFlW5SOt2pD
1UddAlQ6cxQrWg80buLszRc+vQFyqwDtz1zczGTi32QHsRRzsUPJnrTQu3delrnU
lfNhJo1EXRcTbiZiuB84FXb70nGyVdMlt3DJJpPuutoR8Bwaaf+ZDdgLpF6F+Mnc
iU7EvaCHVf/t+g0zPxKTWDJCrMDioOURilKCw89nKrI+51NsZqVoe8TIj6SXcxEK
spjvnpZ+2zVvnCoOl9d7e8ZBPnBXhSd+7RdRou2HVvMam28F4UXqpY7IV0Cl9B17
mGM6Eucki5Ut64EdwKz7b1+BFQdEHc/RovFSC4CXrzfgbcZWcTfeN1d82gXP8t1U
/LMRcWDZC5rjv0y/rt5XVwQkiVr4z3yTqJvZ3NisaJIYqhpjFzg+I8lVQMa7LHD4
FEVFwQPwjct5WKq+TNRqq2YLmIgF7G5FgVsh3x5Viibv1s5JeimdC4CSl2BPk2jD
Fj4fGGQyR6RXaAtt+Z2Jqhc9VHOtOrP6Ocx7oogPSpCVxR2QLQTE1HG+P3ptQmzb
BhDvnvbq59kPVeXXDDue/yIbi9aAO9hVnpmMIsxv4OOqOA8EMmJPu8XCTxC+rpOY
cCXIOgZJIlfTnz8+XyfnXFKiyPVql2EfogE/K0PR/9CKUPW+sOeNMj2oMtijuKCi
/Xf2ME/gwcUgvv99vsLdhZ70ExbfSbWbBEx5WMuMJXiF5Rbb68/xj913PH8etayC
TrmthCTECrAg0mG7gEtK21Samcyz+HrT12wMaHdQtjzCJMQYE3ml6JN6PU+jtn6z
iuDSLF3RH6imWKSphPYaNWz2g8Cv5yMpiOYnmq1GFQHnTzX8mXBvO//xdjFjrPme
+VqKnksMXcZOwjidJbhBzzIc4Gv/ZyuIsxyKMKreRIvmSGT4up1JLcHxP1LfM2Q/
fECQUy+DETPf9J84MMxv6mXC7uBtvG+vZpz9Z+T0jkDjiN3XCwwMvecm1delIgxG
0gmiV/Z3JwIUnu1wUXSLVVMq00thu3ZWBL8GEnvJaXz1jeCb2ktuhRtfI1YOg+2A
t8ydEljYI62pSbEzZPVlQc58aKa68pVZMKYsOlBskyj96gn0EI3bUZQuD6uapjY2
UMZAfCxfeCLAjvPoxCvgQgFQ6Cbyoge1EFmYqRaBoifL7GozzI77JGkWwdPyNKBF
CbFKsKxfShFzzk97a6391bPNNAy+voq0IRwW1e/hcLrkjR6IrZeze/OjfiphAxQs
gINM2z78xRpMJjIvWCyFL6i78urtHLqegsBTZpLQflC9eat85upuLvmO3294bb5L
PNswBJ1DOsSiZK6zAWjyr+KHHDjnpL4pPnY7X2YYgoBzDQOMmztTaVKgAGJek0qN
hwmSboQbhsUWiBtwYAhvHzeDRRdcgl8pHruCrnzAc6kQQq4Y1XPu1rJO3XEIA0R6
zmwLbQff0gOCZLbCTloL7hYpeY87RYMNoi4/B/glFnKClHFR8YaoQq1Tef/33UGF
ovI06fZfcFkVhdHYCxD/jHEF4fW2l9LSVkxJz8iYPa/aOmHM9yyEwO3dF0ZyRhOs
ATdp9oQL/hsWN3D4fK2RShN7KNl6SPFNVaCBztcasjq/E/uaz762t8Np7DQjPIZj
F9dShD0iJQd8uVOXgP+EKEzcykT3qMfHJjVi001JF+tc1ur7vzfO7d/Ff/BzagJu
Ei6Gf3WYSiW9jj0tcD2FgY9Phrjaz2VJOI/Zs7OsI/qpZqzfx7fE+MLLvXek8Xzu
CbVhgUSv679rTl7g4zRNtJH9qIKpSD1Qjm/dXSCOZ6xxgQkQkCt2TucQdDpC9fAi
2R6+2f55hE43Tb5/wwFvzqVk1qb+ND+b/i8BtcPbqTAgv3E8Ml4/PLjkkZWKLGTB
t9+TMM4svDvefsCLAV6B3ARsgpx3rHH52KA24AMW0EXRNr05bpfstgittUx/rzYN
oTx4hd6mgJaHMwU/6pgc2bjuELvL51yjnt5PbHfZgIEDW9CF6KO9xojir+rnepT0
v2pNp5T53pYnO8KZZWWSPe0zDcUMU25vl5BGuS4SS6sftkDTP5WBSNk5vXK86wRC
eN1qjuUCJexHwtmu9Av9e8QvCKu9RKl84+5zxGfCx9M0rZk7Gifl5Da/k4x0D2HG
8Vn04jqdw6ILpOb6YEtT+FYalUo/5ctVqRWcjfm0u5ds7ndpuS27U928YASeXnNH
gfgk2eRnqeYUhJGTpJNwP4RoKiI3fYyTldsuVH3x5powdAy06x0alOikDkIczY2g
BeWvkNjUVYc6PVPVgE0L7pZzbqtJbZFF3FqUK5Tbi6bHiL6ShPAitx28wpi8K2RK
C6aiJx1r47UKKftvd4GgLmG0xCyLXxdl3FROYwnPErRBw68UND4IFyiFNK1yfgVN
CFOduf2h3ibIYVg5kJAmoh35FOQG2ByfZQaa9zyZzggAaM2WKY3EpdDnxzUE2ppf
0S3tlP2IGWqpURWb19zj54/qApYC+tdwvLVzPxAXP8kzCL+kLF2kZ6k2zDsbkhx9
tfZT0fptdh6QHa8YMw0YLNNm47hUwUsyRjafz725vmU3E4HfMV60HTQ38rpDDrSS
lj0NDCOMRof7OSx2uN9wno+VdRxu335oovQUSHpbXjSNGhI6spL9p1xz9frb1xPP
XRvE0fKtif6NqrrVb2yWN3ArHR2FUIY5NCJGrxmluyY4/pZJ35hazXiFtebdU1Tt
RmXfSv1NBm9duHgSrTNgKrm4qrHaCSYt2iVaYqxduxJ5GtSf4EUKnJHj1NMnr+H/
55lUfe3QzBGUTkgAXp1ceV4fPeKJRYAYxvCYIm2cGlPsTinEJoDZuKHNHzRgF/jU
OBgOOCg7nbFM/39zXxWArs3VAsKJPpLAPLikmVNS+ft7OGpF++UaqNyAJ7vAmKKl
CS0EbK2iTgWrG8Hs88ZwhTZx9hzgdro2CDSP68IaREwCXMnDl3pGBA2xE5b6Kn2h
ZNuw6raDEHnInPNwRPuUOvHGFXJOuowVe6cUl0+xDRVG9dry+gvVIhgXvnL+yeca
ihv7WTMWPtjk1c3aI74P/bHAUX+oFZLzZy8SskIiUcrux3Od33As7wRL7otEq5iI
YbIc4o84cv4y9F3h7Ssw/bk72/QWhzyuy49I0C5UBV2e0VB+kCghfGn4gQq75NbT
7jyxFVVZPE5WsOkkrpzqo1fuXSI+EeAJwR5iZY3m7MoUVXN5meAnEyEdSXWdtD8i
u18+t0u/DzF7BQaBVpx9eK0QBKWatzPEqG+JklW43NSd7nNyg5hPxVf3t5cxrEIC
Inzkdl6PCtFEu9ozQ4GyaDQDS9JBkKOau6HAmaqP1XiOg5vG1wcsWFn+2N2dyQtb
iZNCcOK0tmcJPR9ro543S4UGjjIObibh6wrJVpTGjfyuarTI6FUxNleHaP1tqT/m
gX083On/LQ0K1v5VIm05IK53e+AEWRLym5Md9GgW9cWvN+df/WasND43EuC7Qqjp
UhRWkn/sPrR/LzuPhcAfIw+aH+mtVC2NutohQJ6kW0fTxrbX8TctjVorFz5pD8PL
50yZjjTirUklKMUSvyUsYrEBsKAybBt+49Mk2pEXYfR0NSfKQJtkRi0EsA8mZGJB
lpQaOmqEA+0x8iH6Zez1Au4vx/T4B3D+pozj619gR/HpUF7oNwk/4KJFEnLGh7Yr
3+46bNy0hInCJ1pp0EqhY8OUj/Tf68ntIMcHvq0QNwTOuNLfK2TvU9SIKOwrp42h
HACax11bBRMx8tZn6F8TgVkedS28sHz1ZckWJSjY4wO+oc9hwvwl9d+dVb6HYP5n
ABmHBGS6m3OWL7rs4WvcLM3zTD8QtSGQy4IJF4ScO7lHKDmoa5e/fbfKy/nWIn5I
LPCgHNbyj4Zj4p9up33UdJ8Mu3GX0jbGimJYbFNzNR5FChs1uqAlhx3taEn3mcJu
UsJwMliZrt6e8uS3hV/s6MykIFv2ap6Ybn56dnv2GPWnBqrEN3OcmnMJhdXlWza7
LeceYSbTUlRd8c3ICX910msOyERlcsn9YN6OKxwKtZ34PC/0gTkolvPXHJDyEw82
+SGW4C+SIrc/SA7MPygwP2EUhRVDpmt7kjelz3lmGu5tEx0Abnrr10uG4h0XpxLP
N+4fK26yDvQEVQ6oyCoMB6GPiPcuAxLbarYUMTtk/0XIIQlqfOr9l4yBGpFHm+44
oQ3Fr4Hx2OtnR3SNJLJnaDU97kexUUU/RkWTI7qVxVQPtmnRF35/HrnFSeV2WCVw
yqRrEvLXBjalpNiPEsReihkNLpz19G5+MPgOto8HlN68P6wP22MF7zY1IgkUQa7J
cewA5li9kQders0BAf6I5Q9zeWRgW8FCZoROluS9L4g4aT8AQd3V4zC+5HwtOUBS
7I+PtCZNswQegEpgtLE6a6OAOWAobtLuRnINcRxOKlU9cafpWB2Cx8Bsk6bcFlk6
94ZsSTfXv+XaOPk1sXTO4yDRjLy73gPHGD9KNA5I046xnkjLQA3YNbWcsc0K3dMi
/1jwBkEhpXKdCBmmg1OFe0/dyxP13gopQ9qiEFrHXkvROUGf7R4hHEUnmDO4rfKX
mwvgTC1zR8q/pgwW4ar7EilGTGThZm3Vs3exwIqJY8veuxukh2ihcyPz676Hsu/V
w1zeLof86TJ8W57ibU16cScSXfw6hBriUPRFsp8tYJNGdbwxT2E5itVkBY8kjzQ9
VY3N1wqikQgR29WOzm/fST1fIt4kkBBS9tMJlcWbc1mmNXpkbbYXvOhx86EIMWoB
JKIUUxi8ucVlFoYe89v39PeMiyhRYK6D6U7yyMBDG0+jhyw03a6ITUbCqfGfvwDF
OqJblcIS0nHiNrQ3DajDqRiQ5M0j8HQQBdq2CpI1V9uo9cF0CIUfZGGpwgsXOO4X
AHagQqMRB/6f5JgI5kTUNAEhOzMuYAU/noQakD8JPSu4zM/tubu/HSWCTzKImgeL
3CCwHSLKC6/nDaHN/hD9PSHtEAf78bcvW4IDlYTsNtkc3Wy4Wk1zK3y1YTdPvT1n
z/3/L8vSrKam8RDMz+j3A+6xzVMxFxkuIHNnrDfM+TDheYQD2DRZAuwV51ypw6JV
yl75PdwBcrqkvkjthozLAKKHPRgJsN3/DKvjbsMjWTO8PA9z6zxfeixnGXgMPdgV
Ullp7+f47upyfKdDqKNIBxFyoS3ORK+ToAi6wZyLmvn0btj+LWoIxQW60q2T58SM
qTX3datGywiPC+CxKsjOxh7jnMCzF43eiYxbR1UaTNXeW6IqeCm2q72TXhjzVYku
SQDs8JDan8ORWoizA+xaj8oh6tKBd3Dk/f/EVO1hEbr/0qCraKZC3GOln/KmETVp
KkHicjza6geICF+XIYy/he+xogyb2wrQz1C3JjOY20J+hZWubyt27o4258TETb7C
wVQUrrJWD04AHUwg9MSL46p+9YQguQGf9RdKgOEiHnxbKr55L0ew+JbED6wXHszl
6n1Id8e9dS93FW+8+epcc3RlGXVvW2Y4pmUsqsKge2gXHPjlCejWG4CdZrhVCDis
Mra1BcDgBofrwSi6ioRsbbrGHCRq5qsr0w4s6wWc11TqF91642nv0YBszwiSgusc
exnEhUj1W3ctTWC3bdytxxRwITxVl/y+BXCGVPWUfR97um3c1JY32DiCDMrCZbfh
h520jCX9QvzaTA6xr51dvs9uix4p402XYZxVloxvJqGlf6+IkK5B3rs790yBFjyY
0Dgzkocq+KJKav3Rq1y7yBRPIAScVdX/aU5INy8CHtrSeEESXoUDbMj9/CYqtNZh
aCIO4iLiiVvFugrPfddLgWYfgnaL6jk8qejszWnMvwsdN6fFPZ7F8YIP5V1/lbbY
RwFyjDLkXHqm8i7dxloFXCQC5VfwT7MRTFLTcRula/EGOKGpzoJOpm98CBgf/9Bj
S+LvHFFL0+kUVeqJ9l8jdoEbVWAiyKmJiIMmYt2DlRCizaUoezCdbD6LuvdHsLwl
iHCrvwGcBCi86C+L+L3DVobP/vvZ9HyBMMVtYVG64k3tHdNJQSOvJji/D7NDvsLg
QOeKku+szIHJqxTHgQzau+crxR4MxrFzlAEoAj9wIYPG9AVTse6cCuyjYDqfZNSx
akRjuKZgPwkdVU75DdRKWxMMw4EMmfQx2e9b1VZ9oErxJQnB3Ym533n4Lg1n6QUX
mIp4u7hE2Frx71b0KAPmvY1O4a0F9i3T/kmezVy/25f+Ra8i9RhWIPjqwN1q69b0
8k3F+uYCtBTsPIthH/AckN1C99O7xYAg88NHGtyqwIQZMq1pRaajnYgX8DaucMQX
wu+QOsnifAxo6VO2ILkUWVTHtp55xJF/6Is/OjcRxXsic9/M+hHOua9whS+E2Tm+
V1JAlK9/dNwoJ1K6uk3mi1P3KSCMTaoI7X+PGC0nupaXJINuzrnaEXAvsbDeyJG1
uAKB17zX0X92DFdaJRNdUvNt+aLQaMQ7YMWPxlV2aMHhSQ/sSa+T4B2gv3Mqd8gI
VD/zQyK3fQ79XHdF8XQ6W/vh7GE+Zad4d38qVGKrZQ7yv/prXxLXkk6RQBEaF8Tf
6rN5sol8/9rOsLfbuxe/6/4QRQYZv2ZiQcvTRiid4ibCicpyxMMO2G6oZoku8N/i
scHVV4pf7+1UvPXIYFnVXbVinMTbPvgQWrkWH24okLoNmwXhbHR7zDQ9MhcB3i5L
S4z/N8soddv1M1rrK1URBnK/CxU4Yo0OLNFIOJTZ7q/nWyGPhHIniU31EnvTz76x
M1ZFjaQLh88ThQGVSASU98ljIsniRNeSIVmn5sABSQMBqB7oiW2L7txgZXdzXXt+
JrGJfVf+2wB3fmGqYZDzB2ofCS8s99GWOxAqAVRcvbPDoEDvxVJy35ZWKZMh4xuu
g3yCWpllB/a+ltjtfl6J3xHxQMyBKXo4etBtiEm3bcxk5X8Sf8sGITGt+gpR9SS5
335DxNEXIOSOnqCppuTvlv6PdSamv9U0lYyV1aOwjJZnyZkQZMuSteFi1wpsjIif
MIzMaAfPzlj1+DwUPM6T9WRnMT4zZs7oApVm8PdFV9Q83sgT02eTvP6g6daP6HVt
fFx0ZAFDVwfj74utdQO4qqjtBsLkrwUuzWP/Fe2DEJlO707QJGLQHQsNM1AszsUE
jPgA/f+6tlaUT+4gsp+HwsNo8d310PSOf11Ad0Eqm65YVCS+r4ILI3xOems/0pWd
MZ42E1ZZ/SssPHT+QkPFepIVigZ+Dn8FQHpSb2UlywRjGPIt//DSaybUsbzjMZ5A
kv0vnakzzy5FUoQtTxZZSW4xB50see8305TbFTwf161Jxs30jI9inulOUrOMZzM5
/4O/0h5NAi5x+nb4zGKRfLfmWmirKuXo3CXqcBL4DzryIiWzsU6b0XPRYleEyGQP
JIPJKOkf6KJ5PQi/1fRCL1LzUdsZrudzJp8JqGSam2IcMtFMLJEpsd4A+60/NyxJ
acUDgJwGS2EakbLW9NsIwWqRrkSGpYrtuUIApaAGmwj4psMN4SrCatNdEbejSKsz
ZJVe0LJ6+Ikatg2nMSl/ToC2Na/3JlvNGEjsf/0JD4s3fy8VmnAGy/R1WfufEva3
EhCeKsD6VvQCWQuwNcs26K0U4z6MRtoitxNofherMcjsZ7DYTs2pZPEHcpRxrBic
9qixOaARoODkZkFGrZzHZk0F2cN43YE+4462vXMbRDVD3uF1VQVSyzhsXCGZTccp
4M5vvwQEOVfU7qkwVH138r0bAf1HtsIl3CuKJecQzjI/u6z0N6TZt2bsHI2/Ofsp
Pi2eehYkunUNraszN/GdfsBNR1me2mpGIf0sfEsu1dOr8Bn1nDQx/rVbSIXDDos5
5JG/wby/DKS/rqc47UacKM/I4cVZW6aQRFGRlWSMOz+4Ay2AP5eSXRG7v8j6/Vb/
yjXGxcxaj5Y72Ydp/RLk4EBrmNRDxa+NzkxQHvPIIr3bLKQw0yyeYdEsW4JV6wcW
3oqajZA2vRnKUgqxueziJ/W3wXDTUOTfZMeI481jZN1TbLIEYk5eQ5KK2QagYQT/
xiHb5s51IQTLAPbq5sPbqYNX5h1sXENTyxBDWhd9erFwl6/B57VLQlI6z7D2mDA0
/uV/mRMYq1oqH0pwLhLKmiH3Yxbpx2Kk2GcjTnclIQySxAKdxBGhBiwbP6YBDNs/
7+DsCpX3YYNqfqRwjdXORt17jAD7K9SYkN49xWWDcS0dpVMhUkXKFQUVmumXZ/Kf
ICIAvOm06baZkdT5qMjReT8k5kGbRYuMvCnBli/OxsUB3/Woymf7BUXWzdwmicI2
rHUvJPZulfl2FGStm/fHbnyqj824BEmuT1OnE1sb3xksBWmR9SCsah/cUsIK0RPo
1BiMbt3g9tAhMiJ1IwhgyjcKMR1KVi4zl7HGOj6HBIQmzWLVVUKTDwZhQXDarZ3y
iP5V6CQ174P/8mTpe1L82/LIHQQboQblT5FDmdn+JNFSr1oAzc9THNm77v4tW9b1
5w+7SJ7bg4+bRqzvih7WVTl5JE6GQRIU6QNWXj6w22JWbKX3ZM1XEpS9nykecB2T
Mfmdg8s2R7aC5os5aYC2j16BR/7vglTftZrZv4cOcoOAziWrDmxc3NVX8D1u0RjK
8OE8kUowBWoPTkLxRgwLSAphvYXgXtiBO/nvFz5CKsXS9hCptkm/mWvm+eZEVVoo
qbuGRj0NeMQHW8dwOZ0SXuQhfyehDeTdIAypybm8VOyYzYwamBHIm21G4mm5MOr3
8C6Vp23Avqe0fsNWe3ha+OH9+XDEhHIPWPUZOyPvIaMUwq2xJicxktbKPumv56O7
cSgryVN6/UszCx0fQREe8njmb+q2zCjfS6JvugiIBKXra+53QK1CqijhtaRYL35i
D00+f9AVWXsGrPqhIzigCUNGEjYpNrbANbCtL6/Oum9QiLkUPOQcBGDmNGCMK1S2
3EJHh2pbqVB2+oPUA37DgZNvROFkAu6lyknqXFdt5/A0fPKd36ZSazEGLT8tSk9R
Pq7qsOXJ1BdedsAvgsQQ57oaHQQqmWve6B/+MizCiL8EcKPNuPl+Xoj8fIdOocjX
u+JtLK54Mr6BSWXkXG3/+HAlvi1XUJe4Vxr8obE5m55PErFZeT/Bnya2fN0ZoS96
i+FR+e+7BWJACB9RlDj5II4aJN8j/rWfH66TLx9h9f5Ol1KQRvIo6UW93ZWNIL6K
hyIwHWVxsi4cdnxWcJ3fCGZVDZyNNz+iP9Jws46aHxN2UFhC12QxPiqU2tIV6Ahq
pKBQKsrC2xBPvIwOok1TEjHUbvIuhCo/dMDMO1Xsu+e6cbKRtRL93DfBFG3R+f1d
AQV8qVAdY+bn2ecGu6Xg5yI+Cp/mQuryCwl6SQbGq2cTkd4WgqnfX17ZLVQZGtFH
SJdImJqzWo1LBYstrS/UZge2ZFnkRpkuxb//+5sk5r5W7v4ycX0X7VGTai+cZD7F
DnLZk3wTZzEbhad7Vj/7n4CZRYGTYlLYZMdnJPQnBVesPp6Yxg6pZfw0CihDNvHv
W5PFUdWrjIUEhXAw3luIgo277Nnl8NopQN2cwnuvwuP2uA9J4TlosyyVBBrXUyTA
vNYw4vyMWyzXxKhP2zIQ+L0l51go0/zcYJnCDTBMrKEHv2CcDaL2sdNkSZhoDvhv
h7PrDE+Ii5skiQdJyDRlarRSprQeN2n/zkoRmx83IP6/iFX15cCW9NCQ/CA48l4j
enLPzE+J5+pknoTq0aRXNzboOZGRHKHyvlFWsPeHwlucTLrgodH3BfdMTjNkm616
6SJgijMe9wsPKp/tBCSooeIbmes7Lui/V11y1BqJ3Kpa1isWfDx/6TrrjaHZlSxe
yvj8OALXJ+K/dPAwNgAFRvtNv7I8eVKOcacW8J0yOete/cen45sEV1BeP5gdQyKg
xFOLENZ82+CATsnL7FXxMBb42IPvEEbA98i+X0zv2/qh0axCu5QLd0mp+hP17LPq
AcT+ms9RmyXsJuIM9o9EV71pyJiHAUpJK2IRHeanTlunhLitgujduErdcihEaFUF
KtPsDY4apu0FIE12pn3mGiZYFV77JqECQk5K9XeKQ4O1UATgIoZkKtAMYvnMmRRg
V+qo8rgdmDBMkmDdqrIH2Iof9CFSq1Q6IlpVbyOd7xImtU1u2BRRxIJ4TAVwzASN
HKquuMJG2jmbg/S9FvKhknTvsV70o53+J3WPjIawvpGjmAMDgVOKdpRt3oeETELn
pW7a3ORIdhCGNtSrwxHGSSJRer6XBWeMGaPs/WDNdPhbjUr7Yf/YLHaMZSnc1lf0
uSP0mSsTxhyM7YgXuaAZXQBcRoyZCszhY6obHwNtuv5N/ByfrZ3wTrJu2hLOrYtQ
7Nmri2eZ18aOZgO4it64dPd/3vAMWuy1NFS56ZpEsALOXf1DxnXOqNqnF+VVi+dw
j6Bz1Hq/XmZ2WgXc43Hg/PRFCc8/OJUBxjb73bs+LRlpRjLnlVkpRBSQayr3cGUw
WekvvGpXXPddB4d1zmXeuWDTnfqY+1CDcxPPKxRnq6RMtHtJcx6JyRsRfIL3MPNF
GwB/nqZ9ySMeheCuzM55YV1Xo15OC1SAiP6d4qjmIS9L8znnputiDQXMBuTu+J+t
K0nlg15rDoAgDsv4PLlfF26k69EK2BG6QYnfWu84AH81xC/FMsKCQbJwinrsOQHq
Qvb29+7jGtWS37TSX3JXFXrT/q8olZswrqvZQdTY6GyRzQfn75nTWe+hY3KhUVR1
GGA6B08gEHa/9qDtK0Juu0pGOMo4Pw0T79RYYKSLj01VTe6wVtrOr+2G+ZQVicL0
rJKwwfUqgy++a2OLDsEotYbfNrDw04GwgL/FQK+NLFLXikReGLQcNVZCK2jiQYsx
z9XA/oy2W4Xk8no01FawTjElLen/H/C+i4dj/HlIieO2B3MFd47QFRCgvd3V127Z
X5kYEyzrg16yupL1d0S3PVDDqC6+uqUCbiU/YVPTU6uEFDV5ebLLwvVm1zfkebYe
DoIt9bE6QnHTuGVKjYBLzLLKNMPAbp4xMa/EUtFDGzo/SrEMY4hPkRaLizobGzJ6
/LqlexdYbgNv4IceKXTd8LTahWusEZFOMNhru6GSTMDlh6hbm1toT/NUKO8nMe91
YwCBnNvoBfi5j1YI8IQBe7pwMrZecVz/ouTw0IHR48snIE0Obroe4we+Su+ulA/2
5DtAWiFVh9E9OQWps35yzIKJWBOrsMwwpVOFH3KvJJEjqKAeodvHybr6KTzVQUUC
OCeDHvL2apEeIq+Q2swpf8ShD+yN1UOGTIqbp95nr0coyWd4aNFNXRRx94bM76ca
Bk/9BdzIi8vsJYCIo7H7JXMV8Uh8Zq0btbBAZMBkVoTLCoLIni0AdDSnYd9phPhz
Vp3ShICwgmDfs3EQVFQSBLD1ZxDDSoILetJV74SLuSB0LlnWg9A1noXeoQOiV88a
gRhgdDg0PKZoaNAEOw06tvt/9TWiTRA4l7HWoJevf4/6JvHMjtHwr4IlOWKb4GJS
SdRtdgEvoHnuWSzvEmTfiHKhEV4XJ5QBUapXMhhgzumrYvwyLSWrT1DlSOlKoRNB
FGRJKfhRejSmzKOdWFEJh8qMMasGBVnqRjC27jNBuKvMtmm849IZhmz+FhFTyejt
967Auhg/Z8mtnGgMHW5aZjTJW4mg8XjMbrTSYqZ/Sl+M8SZlY9WWQUF94eIiT7wc
n9el7dJxqsn1Iik6yg/OuukRArgRXjAYfVbbFXslPStc/gc0DUEtyEWGuE9loZcm
Nl7LVx95fbjoJbnjvJ6JTwm8XlmTnV3iR5649BnuOFD7yPNRKs5pyfWjvC1Q31zA
JsR1FbIkRRlhAcvk2mMUZD/bbRJTIbU24umeWyeW0UaceTA1NOVYTkweLgqA0Sg0
REYMShbTh2tQvD/GukEGXEB4v1zrzdFECZJLHAD/bZSovgGOVFvpT8eVWqTAN8mV
G5nUuLvYyJ+UNP1F/86mTaGB+QfnEZsmA2G1aAnNSkTlwMISzE0MsXzBpjCk6pHl
hpwB4CfvEZEFjYgSc+QYk0/RrBn/6vX3X6SNPd7+ui90Yjk9X8dG4j/E7KAHWG92
WnSPpCC1Jniao3O4HbQwXHtZmaR7CtnfegmfdxqovWuoq2LVWFUxUs2lskIWmoXK
AgvEDrCDWkFhmzOqoZNJsf828h4Xkp+B97MWR4f+PTFxB5NOS6om0qfR88fW8GTA
k2fHBGLz+qQbgVtIFxNKKgnEuNyXFdoWbf1x0c4oXRNjyPV3jg8g+D/S662cFRXM
wnLYeoZ58VCpAaz7BrVaQ/c/N0E9MDOlQEqouhGssj5a3P9NALTo6efkmnoFESjs
4PWcBxQUF4xvcife3zH2sWpz/5vJJ5R5wajQntiP1fSKZmWffTa6EuMIjOdMgfXB
2qEMAFTeP5HAK4rl1i3ncgX9LxM6q2jLrT8W5g8Uyvf8tHHHtRxrI6Xy64TXNaEQ
XAe1SybCrRKsRkEay7cn0yQqEhAIjKPIntD+VJ/AN5+GnDxA4vHfwxwPhA45pQ4k
PT9xRsi5+UpTj/5JkRGLVNYVqwyNu2+08tm4flfnT2lN5iZjyCiBRdHfJXppyFCv
4pyzsoiU7WDeEwTCQ9LUvRn1x4DPkgw4QP1y7uHXcl+umImLjYXUifbFG4AV7VE6
sA5VmIbX1Zl90IQlAFSG/jDH1zDiPvtulko4E16r/xPjr0YO+4DcZjBeFaq4sWdx
sy+8iPmn7CROpInEgx0aPmkp3RBchzdDRffsVtaDI4HcAg8N/NHBWOMadovwT/vh
zKmGAgh9sG2IheL67nWgVE5b2oEQyoAqSYIVjzR5E0dtC5rYKCfWLHCab+4jRq/4
0n3E9zRso+fEt8znnDnPHoiPuyHpg6P/CxSl950mNyrvMZ5Lnfj6OOY8/pAbn+NK
VQS1vG9DWyJ05XmX+sq9m03kBkfWQxE8yccMfrXv4v5rihL21XBebPXfsVW/58CH
jdyNuJDgucomc5NiePjgRvmdnD3OU5KOqrZYrIpcSnGaU1/ixtTlXmYGbyAttArJ
vfDFDPRZcCJ55gwF0HpoeV6iJfxzcfajnjngPw5pAG9kZZXsFUAMMvtt9gemtNTh
PfE/5cA3ihn8bYkxylKRhczY3QFo93fqsya/yVW1IT8ZlNiEfb8wq+XNVCaS65pi
0BD+LsEsE9gW+QOd9r/QQx65n0oN9Z60LWWbuKsGwhTnkP5da/5pbfrquV1ljSV2
TedTmk6dNEOSlU5yCp8R0C1ezS1u/Be/RgPYdy4XZtUpncbRrf7Moa/S4hZ+1piT
RzvAUE2m6LSY9/KYIu085veYTaTJW/vS7S/s2CAmifQ+xBI5W2w82QCPYeQp8Am+
HbvQmpjZmVRmM/sGY84azkMGc7YxHF/ELaq/9izhkrSo/17nN6zPuuk7hPLxpHgC
MhdJnLL13m8qrIjT9pQyI0+PQjN5Fm3Ii3rc6tOn56X/1gQxC+SFpA0kLXvGGZfE
iMGytoNLreWnHprwsLt/eLSs1KMlUqvpDe2hU/egiOXXxctenFhaU302yvRJt3Tw
9Zue6n6MbOZuAEYwmuL0IUDY2zdoZhcqaKVzyzKjWy7Zdv9l0fQCf0pVkLU3WSbj
iqCUrm0H0tdyIx9Y3qO9nkyHOySFxD5p7SSJtN1IIIK9j66qN+146CMzNIueQ2ky
lnKFymKklMGu9tXGJW2BN94wCAv3b/XM7d88Z1nbz32bsvinipuvfmQ+Cb5SnwXS
RAQS0EVUMsaiy9PMuEkTbtWzJfyG7XovtseAbcqC+sVCyDlXbeGcWQf79ASIy6li
LwMq6lZTQVpqSMuxFjYazZrTQQjpe9YrO5MfAtFY5V5ih2IW7zpv2HxmEyU5N7f0
XsaTq1LFzZVWLDcA9ElkXSAKcm7ssG2pspzZxmLDmPeYkApkaUp18cjUUA7uOEoq
Dg+N1VIvSuNjiyM2KwanXw6Lt5N5iXlQoynrxE0JHPTW4iTq4j8yUQnyMtXG/2Nh
GWvc4EUZVXdr//CDoDuxjIuT2hxt8Ln76eRGctJEMmEB48Nj1uqrDfjJLzSJNfG5
OUJUmA8MyBqd3NYbo7ucss381sUHWYJd8BAYckdSH3IQ6+0Y5UBp5TcIuCgYAPMV
jIdvFHz84Yr3rsAo5hZyIQXr18TyWxVbl7jNqyrUSNVrOWPjFHq4PwnoDgJaowwv
4CHulyF+yIS8oLnepMzzVNJNsBBCCO/b7BupDMhI5dcBlLcq6CcIiEDAzMEVmIn5
nmzy+A3y8wng6sv5sEJj/OT3YKoTfqzwWkhzxcCX3dOprj0bn3kdNNwWokZd2Z8o
/2pjARDK7JctWZtx5kWmpbkItWeGZ1+KivWLRgwkYnPOjB5qCdEKA3Hr+0zmFrGo
X8oMyPY6OV/uFbZVGUVYNquatY0otVM4FntPGnhmWfRsBAg5c8l3AiP4sg8+AhkP
IQjJc2NP3if8fvnrZHkcQnRiLTWYlMdES1JSfiUs0eOGZrgV68N0dE4YxDeIPF7t
QL9cAvNfIZRov1yxfV6XRi0Pu2Tkls6bK8aJNfa9kmBZ70Hd3qh0EmXUTT8am5G5
vQfdKf+UzTb3MPz2SEmyqLnbzRnLsF4bbWk9sgPBIR47qwKMkFnVg+FAYvsOTp2f
fkt/DSxPu23+6+a6ax52JpNGzPRew2Nc6MeNMnbVnr2eUZLutmDh6cmwPTFU/gMg
Ku3e3PNveDESpobVL/PerFQwRd6h4hRJK5FPi83wPXZP+VwQ3ehVrnAdg7vi+xLZ
EW16XVceltMdB3DAFXSMQ3augqub0FCKJuFptCwgPeUA8FUUpjrsoQ/QS3reW3y/
4+KZjtu9Dkt+13rRJgfGlYZeYDAhqOOsvgKY5OJXMYWr3VsFiO2AvkWVRpbxtnbs
J2Uhv5vlp0ubIIGv6cnfIuquSehBV1H8s663TNlqIQaj2u9gO4fxlhe5DWzHLfUd
UBbmZRRyJUV8sl6RBrrFhod9C8Bi1lnGEZtEpfgKrr05a0UcfNYsGzbVDtqszn25
1M33wvWs7HJzQdsu7KNIxrHzKbICytrdDCK9DELnLQhBPulC2Ln9GlC45YUe4fhB
XIGmXQmV82Yw9kP4P9kLutIN7/Y1e7ImvunnLiqQDCq/fBeg1U1SWyPrBhOlOZC3
iU5G0Db/RN0fv5aaq2zS7AzboI+v53YG4P4FTmLrN0+45yzwMmjE9UHqEpT1wBgw
bjF67CTIWxj5uluIwjVWw3Yqwj37aiSOo3EkgtZthrfEyPXy0qG2MEuEjAZENUR5
+yQ3dmj4KJUII7+cNCGBZrfKSm+LjELL5RHP2VfSBQicMaxzSEPKrmeNqJaf3FwY
0r8e6EI3EGVTtiTju8DL8Yt0aw0k+iUsDRS1KKotN8Vc2Qr9PvnbGjXytCXU/Cu2
OgZ3uWVixHzlVn/vrabhDGvbfgUqQBDwDR3WE95vlOjsbxTHLgDGEQ4ymwRWJHx8
2PgjIUrY5M7v3WBLY+qqkO8d6y3FRyGvVvMAKMOuZzhQQIdLfrIwlacSD6rO9hJp
HWfFIzbSFQILQvr07q1a9gm49N4DFdCZ9rp8YSHnmMIBzLhMDz8PwVdqAZPct2OX
jWZQbE/tpottrZC+nJXlUa+nOPhnc27JOP+fNQv8HbXXXZp4RQ/e+uqrqRvnnxPI
Lw9aUGFPTRdsGDY56xaiHDM/qIdKNtv/Z68tMSTU6K6b7/RDLLs/wV8j6duRPCcP
uTzfYmShft6fcwZ99Ur3IJZHx+wm90aJVLXN9ihhUNdCz8q8iaUPTtwFYlfjhztw
Gj2x+YzV6ZnufFgDeQDyivpEm23bLsHMYfQ7dyPG2wYCVeTGsq38YECl6qURrhd1
OzCleKq2kkswjy8ExtArNwoStxtOHh+WF8zdFx2JNOKwiC2Kav7vIHormdBZGmHX
w+CRotfGz2lTYxpTEt9XWkc7Qnp8Esddsaa3l77Bla2R4pGowhTi1nxoHakhKs4C
GldpD1jdDJCb1RlipP4At5AS3BmZmFZXRMl2xOgkZwxDC0XEu5Aqjvkjo9vIg4jd
r+xJqFYMwxIHe0ThGvAQQ7P0m4uWiaXqTAk0f/hfJc2m0vuSXii5FkM2vuzu5t7P
C+jvGLYOty4OguyS1Y/XsedD3X3nDyOIxyxybVZz1/gMuyTyMPYBM5zhDHFK5H2O
pv5DZjOxn2DWjzczJrw5ZjJFjC/4XhaIOTZNG2zQtiGEl72gLaKZV8JV9gQF/qMm
CtG8EzDKgYO2gU9TbGrtKKNTglbJzJvNmnoe0ZGKNns3OMbJdFyzwYhVFeijS0Di
L1dCHbpREGbwWS0zY+acNieNAtTLB5U43qurla9UzxFzmxRz+1E6zJDtzU2FR+2o
Bp2jdeuFDg/+Hkt7Qzm0TlOEXdQuqeZ9g8v915aJKVDv85iyCjbyxOGRNXd6y1XB
x/ShFRjFizcseRwbs9e0rosCAlYR8jf9754cYyAt+G7j8leS7a7b6VDRYgkYpksb
0mUfrRTLYmFj9n89mHv9/sTHelt9AI9OGI/f4Plr1acEfHNrmVQAh+P5QSvWHW9O
Rs5lb5vh8xg8kruoIgQJ5u+Xg8DFZtgHn8maWhI54O1CTN/7w7p3xBSI492U0BCx
4rlJTL5dczoG9YOazoB6RN1wedxHXQOOOEZjOXXItMv/+Vu8DvXKGGQ+gKu1Ntzg
kNoSs0rOJm/qbHX7ipTOvVKwS1otbEL3Zmc3HQfPH+Bz7RVurc6JfGR4O9iG0f2W
9Vy9kz/TVi3H8CBGg9xISjVwZuvMs6tobMLuNHPaAIiUUEydOERumKDB7YM5S6In
70R/AEA7TwTKtM4ttsPWSZrJh9GW23GTNNc92dXwQ61f4qNNvULWla2cbBr5YGXb
HZaxU77pow8JB8OvfKlNEt89hqFlwERoVdPuPg+BOerQK+CbKEhq0/yeEuo+c2r5
/BldgIWIILuGfNxqNpeQDm7AL/vUSzZ3wfhWO25QUb7aZwh6zNcmpAgewPNugQMT
WpH3Im7bOV914/CwoCwWL/USOZl5eOzyyFyb3KU3KuL1hHVnrQDMGXe7Q9fnhYh7
QICI3nLPXiS5wd7EFVne9ck3hGrEzPNSSwkVP38zqyFg1gb1JiNMcjZCxxC7MBQ8
BhutAs/Ux8ECjJP5lGu9mS3wGGnwDTKnyOCppVPclH0J1dQK76YhnPgnnbRYI4Hg
eITpaHwPjmlXGn4dQwptDmtDSso+0lDwlkPTbFq9MP6JKM5v8i41MkIqOMwnHTTv
D/Cv3/omfC7+aNba7BwdrpLzO0rd0miJDsGHylvLj6WGUtwuS4kBI+FTV9Yb4Q7G
a7WRm90fU+8bqmuaGrPfJxIwn7QP0h+bGw3AoDMuDw6Llarr02R0wCTY2j6W1Z0M
O4pvAvrqhH7FBoyAMokAyA9TTmxlRQhFAk1e9RMjRy5htpbwLLJJxNDWH7tnZdNH
hRKZJgMpZMwTifMwItUBOYzQOuxhbBeouQciynSY4IjCI+XwFqMYzdlkflj3Pi4k
B6KAihhFgynHaBb+NMrbFgyjYy3qokkU43e82XYs/30qvkAt47QzRzxmbu/Wlqqu
5fGj5SD6jKfTZq487SP9bL5zJiAYCjfSG2Q4x+FAcSl4CeAowBP7HeH4iE3QSQvF
8yH4NTo2ofdUD1iLsccQa69ReU+Un6vTjpn3Ad30ixLNZM1Zsaw8buf6+SYSsN/g
kePYb1/KD0cPy1cjljGQAVZHAoP58ukVsjVdTlyJJyE2nJmxZv7KDsVbfXoB3XLU
xKm8J0mp9Y39c+XsMGoBET1NZPdfenb/95doMt/N1qqJ9pBBpCYcgIqOKpPthHhn
dCupG0S4ZT0nCXb+Pv9HZUtF5mGGA85eH6Tv2tLZjO4XoP/C1ZsjyZyGp3JsaxgG
Oqf/blhyQwj3/sq5T0Hbtph7WB87agMZ+HRFAV/ZnGnReW6OCYpzuOwaoGF4hHuq
Z0YDa6XEx7B5hwh1BKDCAEGJlWGaLo4VhfTksDk5qPYzK+q+Jj2d3bpxYaORqG/E
9gZuGPzPSDAbsbTeIT30X/HbHulBxrdUKZyQFG/m3ttvJM05SbKrkCBTMijH4wWG
5BvpyEpb3fP/2qojWoKHOUlUKftI1qB2+TuDp+n9yTJz2Lig5mwc6sTto9HUNRgG
SbpZ1JsqzqwnDpakaNPhRhw8HqUrj+Rg2cZKj51QsTHGSxhGvd7CdzF0V0UsZm8U
JpA9PlV/cLwSpyiVhAAQlZMLn8wF85Yg1pQrTSUr+ftIUM/rSGdaG30qtvJnX3mE
BSDQirwrGY0dmHYt6ScUNO/uXy5agWsxTSb48jC5lnWEVh4MyonlQUg1o8V7x7cl
NBqNK/y4wtOEdg/FLn3AU5KqC/MOI2SdWSF2yf1jI+7RO1p4b7HFWMYHLThfsgHd
extYhSOSHfTXteOS+JBgZPgtDz7K41CyCDSdHL3/Xs/Nwj3nUCI1STEN/S2vuopm
YBHkWQbG7WyPllt/J8YJzrdoIhz0iTXIBIBNA+oEKfPoF/7cP7pcnPkWtqywsSI2
IrvrtEN1XwyZL7EIgqme0p8Jnl0XdcsIZHlFvflGH0BJsbk5eVtlmC6+SZpMKIsM
mRcVcY6dyiajKT8CS3OhL7bH6eEqnSU6jhjdm0OG86KomncvCfjtPYhX2fW87vQo
deGt1LdPVlEKPDh7rC3o32dJWWTo0VoYr7GFPqO4ZyXGdRl6fSTXn9hJaP2ZvuDn
INeNQbBc06IILopB3r9NPM2+Lano1kME2lC+D3x8z393ub2gri4o/0Mgu7Lfvf7c
MPQ6EyF+UMwO6lBgwAd6ij2z6WvuERWFeJ30fSyIysPGtUmaNrfYBJVWzbTKnyw+
9exfc+Iwhw0zAzKHUsYGiiq81AP0Q77exAYythgmbRRC9TYwZ4t/jRf+OokpLq9v
bYCWfZeDQBC7yxUYi0mLXE0fxGLKVM4K+pP0+U1N/Cq/baTPFJWxoulPjRu0z3s2
8vtq0yGHQ08RBDtLhp4odCAWX729nBxCA1UXpgtyU4+WUvMWrI6JA4WxUz/UWJBp
rW6ILexj2flPRYAsXJKj+PuWYImV/SBMHFLHCaUh5+BoFDOZHUYeBmI16ls01Tw9
RCXcLuWc4nIlVGuRZ8HsOB0uAiOxIMP4091azNBBSgjzBJds2DL8e1Elvlj1TLZV
f1yb4l+mj007PhBUNB/CVlS/IGkgwGdb5XpDd63ZwhVtIsvo4xQDbPYSHzwS6u+/
fJKRjR75EkO0V8GfScTP+vEu+avHCvsgtlgMILkMFRBWi0BDD5ieyuw3XwHoIdnS
56QoiBvngW3b03B7LNMHnT6+kDYdAJThaH15P8jXGKX8FK0BFgqBhrwSJBIWbR4u
X4UKxZHN7P7rsBXzjM1HEU60AExz8l9Q9QhtRdvYPFv3ifs/2U3iFcrbCm8qkBDF
Qlt4pEQMcnkrOzcVJ3I9ScmCyoWb0IUVvjdVMBc/JsWW0zJEd5s0wR5nQ+HRk2FC
CBumidz+2nM+HIG6x+AAm8wQ2ahf80OtFP2QMN3F9CECcn832kVF8wh2+cHq0BNs
CRmbh+uWRJ8h8LMd53hq5sPBSIGJk5LdYfjWBMmb87ltQPk7UzBJOEKFZBNTBd6z
3Hjw6j29cqzxRpRiU7yJDMVm0ee59PHYAnVbJJruZMifEi4msk3jjvUnd4/YtggJ
I4nAfEjMQwFIAkNxHG0zq5zI5hA5VXFuroVAGldUKAkhUflqX3mVUVdjeQAFKiev
cFG2iVniVZbWOhSLp3PkVQFH6l9mcV7hWHsZGuaSvSWQEFYxwMJEhvQhgV/6Rw6U
k12+ybUdfi5Y39zzOot39nDEf+u47i53PDvqzpYFrFZYX1wITKJ5FW1dA27mOqg0
RN8Pjg38AE9P81T+d7lsOirlZ58XlQsHC5TcQ5aqomJhELfNQAJxInlbdgiuGzYA
HXRFJ587lMjJbCLijqjDUjFfnS2aD+1MrQEsElXd2YqNZhb4BYJ0y2UUzYyaI4o9
vWzcmdq6tmlEXWXf211xOkuD+h3I9mn2bUbb4Fum7au27j1FyjjMNYodjzHe7MDn
NgdiUUvk9dzR9EBvLJHRSXrURj6Hz+XnUt1oHdJEoufyTThqFj83pCtCp2ioBF2c
6g1eoCZhzjfaLiC8oSBVlBwm7diB/X+N8J/C72q38Jh+W39aUzKXXd5MynBkzQwq
q3V8H9fZOZvGbZmtopA2BdDKr7Lk9glw9MboZw4amTo8lcDo5N+C5vzxkAT98EP2
s2kvSboBzJCA0PYEw1NGwZVvKE8u/NjGH9X5DKjw7G5iYvOTW9VufA/HCAEJWHmP
eluO5IgbQnr6O6aWMH8Fve7rnXtUv7qpoae/NAKCz5+x22gEGRNBCSlzq35cZubx
qoI8H/qd9TZ7NlLBZnSX/jhquM8IaiIM4CIB8NgzZ86BzVFmq/Out94qAD7LMCRa
HsuA0QATKeWUYwq5xAw7WDno0hlQvp3cNsDV+QO+Zxbb+RvP7CKZEltukLGM0gl6
vZDg6rjyK2h/aAZzHVBuPIcdyChXloIfbKVARAoXC6Vz8/Cd/OlAfNFpN/3Bnqux
PGDQQ4IWaCX73ysrR+6fhhHmf3qLnjTzM1ksKaJ6CwCFwb6Gy+SKXk7Zepsw4UYr
McBH6tLmJc+QSF7HGA64mkidlN9ggvg1oy+71stB9WCqNzmnjE5+e3jkK7ytg6QB
2Tm3XYxlTvSUDVGRtuNqLmPvmHiPOtgz6Re1zVLiByoNzfrCBCa2bLnx+IZlW8zp
0bGip56Nn0Y+xlBbW7cxfQ0E1M1TnEQrgWuk4Yo9pmojg/sDaKShkp03Q3gf8oJC
+Uu5/PkJJEqM2TiXFdB/bJEYkfJpaX5pEzNYOEaTsx6U1gACxG73PvuSMLn2wsdl
AG3gm4rkhAp6YLS98XwPlmGptAulhMXyNEZBuaZKNg8shpmowxc3ttqTgDmpJSE+
JapQpHFrVAalFqOZVzZU89YNKVEgneRUuV09PFtYBTCjEZYaj/UlcP60u3VLF68r
tYhOGsa6eoti013rot29HITISeG92VQ9vRJAJFUFsgvNILYxcoJQhDVNwh837ZoH
vPvdFsdVmQEwVQ5BvgGzM2eJWu8S9Z51Y9Ol4iuLEbq916TqrJZv/8K1r6IwzXxP
x5LtYDd3ClkaIby0FcD5mb+2wvVV/iAEmHr/Ngk+01xzNkA2uM2TKrtVbHLXajd0
zap9EFJvEUIbSUlFjnfUuxHBHhT077h9QqGkylirv2t4iLTHOOmR3D2ZuyukC2C8
NH8AseoKKufaNhqwfQGPlJWfqyb85MkmSSPFfPLNuZuYy5GhyBdQtEtXwfTXdTIE
sFjN8Q0h7nABuCUHeSiNeV3QC0sYEYOKG78mrzwlJY5VEkcyxdXpkLmwRSfOnhHN
i3+EJSSm1b5buh+OlUjSw/U7hG3Hqwszd5gNTDEnLxtzhgFZv8Z7ucHPJ21xeLgC
FdlgGbIcQP5S+I4gziX+Gxu88nS617cqfIVSJdj4rYA3T+6jd6uUDCd3OtfDrwYd
DJC2rEOdE69csI6GYxR92/nxi76eULZTk0BjQ8waqw+YWByXPJWc+Ch3lWd6GpmG
Vx+/1rCRgGE3xThuGL32bM3TViHDB6tYkGYA4EmOXuDEhpQqAbOqXHpN9FktUasa
EgLrctdVIazVk/P1iUIAb43RJNBvUnLIzfZHN2kwl8a4enX5bhNXkhQN6tNH7Jhg
4NQRSJfZQp6imqBmbEmD8RrhB08D3aGHeYjVKEI/68tLKN+udsy99fU/l1YOxcac
G+Wl0lTRLjVuwdD5KqNwzOSsEBx4DmMNgr8ylPvx7BzPpJsKLGb2g1xqIA7af9+T
0EM0Lu9caWEY88BwW2gN507BN0MI4UpK8/B6/6h3bwzQehxYK5vKr3bbWV8CEAAu
KfUBqcUvupZMqfwmplAvuz/9vEFI4e4SSRQpn/1aUcHpBESNywdj4Q7VLGgXnwVT
WtjaHtOY7LHN/uXBYRRXKq7TMguZATU9y33qoHTfmYrMG5xUwNFBPW6E4Grxayoh
RrIbFPUbd5SB5p5K8NRSvoF4EAxfBBsC6R8Lav5R15T2izkFaIZpPwys/6KbYBAk
JTXQ4SwVv2toeKWvBaoO9wINUmK/7LbThN/9oHNJcWXbTJQrSSHlBGW/gj367zdQ
tSo1x+2nnXBF+fTJ1aU02DIRaIH7RWG26mP3j7GbJorQunDa2/2E52n9FNSxJ0Mh
fd3Lrn0kT7/k/m23fJj0DdRFRcpCXwd2U53zs49VFX0iiI3YW96ZOTCIFQMZU6te
pLN5Nti9Iidh4arPE99+5fBZME+LMNLUTMNGjHjeCFiAYLjJPvgZXz4qP6Uc3pxt
Id8xcGiJCy3Ea5dmBkt+eFPDZ88KRCQUDNNoutEJBNTV+hnO4rFnRemAiX8aPrpw
vbVhahw9WhV1iUPlf6BQBjugZd6fEpC1naNtshEye8ybSuXtUh1RsiljMMhCG8P3
ollkRC9rxWhep9EFThjCscecAXrYF/wxmdKmt8h8Xgbu6xKKyUaDlRPqtrK0nyLZ
c7JNGLKAYP/BlPjhoPdaEM7yBNIzf+8hYQja2pVQskIaDKbsHTbw2IL/Uq+piMkb
xBg40CPR0VlpgRyR8s/dCCYbso/BY7jrQBjk7ROnf8q0JT/ntlOBvlzJ3SF0fp2J
roxHfMNhoE695dp7LY32flFI+sM7CUE8/0FIcYLGfnSpWtsqJyjYuvHyZGz2JSMJ
9hdkqN2nL1KlC1JJc0z8fe6a851vWcp4Mt2m1gpM+p1mFKI6XPTZNbwFUUOXO+WS
XFtsTYNPgfh2/DF/AoIuYslCFIAi9ka8lUfoIeUbMV4C8gPASr+Dx0wTWRSlnHQ7
GOCic8jPVBsv9c5IrGNv5cWQOAHwT3VMyqI9PPz5S6PynqXrAmFi6Sc9VLr92+Zy
SZHAvD3D654z/MUOzouc/0rDWs6kX7LmTWTOFjH2KRPFlXatQq6frhRC66Dy8olu
eOvqpBKW3oztJ3xx7S2NNBIQ2WhUukBBVQWawSfBKekcQjulQmHSKFx+dUGxyrR0
jyMdTZRTX8yt/1f5211YGkvx+JImzufvKCiJzQBu/TOXcmi839uiH0V82DGI4pd2
dNUqhbrsWnoVH0iGmZIGZqdtrzTaXr/SewfTo/sJoJQuGYiq2X6wSssQLvwY1O3A
vd1BlfNdsVuvnrRY6XDB+pNlT84A1F1QtVh5jctGH+j7bXBg01qjLabsvr08knbV
rTgxZ5MMiGUplwp5L2thJhjbjrmew5UEkWlHy3nPJpLBrYg28/S3mmN+9dfF1EZy
labAxzKbzrb7beVjxobb+v16p2a88BjcOZ4gsWiffbUcxT3VTp37AEzfy3W3B9GX
rjMDIMhwkXvii7InidGsCKsRUaOYuQzgqQWgoMUKWPmYs4QqLCpLeRlTbiG4NKC1
u89dnlRr+y8BK5umAA43uyLPEvnC6KlhHGrb8FDVERVaWfRFhIx8xARj+GbqPLQi
zyqSIKoKSbMH4GElu59DMVExjoJm44kzYRfVFMJErO0QJH5OoWwA5uD2kNQ+Y0Tk
Vj48PDxtXXjjUAamJ075tP9gbIfupNYvHLCE8d2Tp0HMNe1ulbNu/sjfqGuOeC7q
2AcqfBLeK8jvzOVx2dlHg1Nhb4IwoOdngXTxYr6aHMvRFae0m+eb2jDB/RzqZgNp
aZhu0YvusirS98h9dNv/jKKJo/+yKnvSlov2k0868Fsnvg7CAL8jG7orjlJYlnMD
QiJk52Ev6DVvWOYiznQffV2ZUCCpX5OfdhUyA4iNDKjZQmf1K49twMz1berGjUvz
HNXIKHrROhdMWTD1IrFy4pyRmNQLtfAqP7tmwHlA9MHgGMXvWwsc8N7wJ711KC6t
mGa9Xf4IPNaGmqm2lg8SCH8hEKGKFbgpkIrvh4fQlBxODWkhCUgBzgf7vXsX89QX
OpEh1etgOQqmfIs3W6yHXfWXWibLkCc15zAnUd+uITrUmYRzS6LZ+zohkEmYMRUX
b2czfzi9Y95Hsks65MoFEneQKh9dgM1Ck5axiaWr8IX112AxO7Y8G/m4MFvFc6Ur
hqcidwNxRnZnWZvTWeUaTd0VFaDrbRGzhXZmyfh3TQqgNwHxaHRV1DboHt0Q9Gjf
aDHSPYVDXIMGKba0tfK1FBdmg1Z07UvxjtUy2jwwCUq5SxSfkzjtJPcz6s++bAJ2
UGZpTPsxng1P4ZVQDMVWBN9i4OQ86YgNp8LdIwO1sRkpBoydUnaJURH5LJr4IG9T
RdTx58Y6B+XMjdlskLLiQJAx15v+9ZxvVm2Eqqn5PXBkMC8dSIPnUm0OGgJG/EsI
oxHHmXo1t+T2NXXkZug0roVX9s0DigS2tS/C73DDkFRyllJ60pUhkpeofiU4iLcr
6Qe6sp6VRYO7EA0vnElrLcbesGuWswLLBeXyHH0Cc8NwCDqw6M4tgULPh6pR8fGM
byvCaZRLrWoPMK2z6gOloUuA1STwJmRMowe8X1xrgdIGtROb4GAA1L/hGNfaAgAm
W6f/R/0oAIsXNcUfddpslT/aI+CZy40ajsQ/OJFdadVCf4+CdF7UMPUlgDJoWCzg
v8qZtYLvoAWxHsZQi7KjBYg6HnM5+gyUD+Rb1cQC6jYu39xOX89EhSSIyIdYCj2U
zIhlp50k38F77Gtr4bIyB9p/sYPHERulduSgQzBeWS1dJtT0ND4CJvelQYD3IXzo
kO6niuj89ydCODLxBchJPPqqjE/LUBc7TuxElWebwriVW2Q8vjTACr3MXpdEPt6x
ykrhtLhKb1jKEOiT2fpVvIxlPVhvTubRauPk6RB/VnSmsJ0PnctCdHrUPX8Ihw/I
bBMFA/W2hZ+LbJkQBeIlEu3dh2AP1bMyTXya9n3lmdctaFTefHu9tiXYaSkaukY2
kpIHrDpv40rBL5MP1ok398OVKBeddDB8hVbWgiMeBj5qQ9sC9bxlaD5gk7Bdd+YL
qrBqBwZQQDXvwiEXMA124njqzJMkE3YzZTHNRrkGNo2r+Rc0Ey7O3bPZB3WJXjRp
QSXiK6nSB24QDMIjkF1LpBlYpo1QisWOSqibVDd/8CeaG8pLIOmJgJynTmq+jz5p
N3fgrcR3qrVzqUsgeP8UdsOdrz0dPD8kXmuSBR1iWsqpF5aU78e/Uiq93FQU6o+e
/Gm1M+WcuqZLlJ26Nl1i5EfahumKk+SvKZVocE2VRFgpLMJzM7l4vk/SBlL0Dh66
bvmRiE6x3cpcUzcX3J8ZMRrhw7yW6X/DIbyfFTP7a8cBAuePMnR2eHJXRQmXQBMB
rcg9VQIw+WDjhvXMUoyOV535F8g86InAuLl3np8O4jYwXkaoNfqyeI+nIvl6M3tK
2pDxFFUBzlJXmdfnxcRPBvdqAEiEP00wPjFCo9eT0Gm64CVqknP4Blcb2ZBHjTVY
6WWVM7xSCptxn/N3JLIYj2o9bwz68cmKIig5c0IotptC4MlrITvSL4UnMCtXMuUj
jsABBfX7DRqt5N2jkbe4tM9+TCd9UWTGivMS0xcNGttm9glvLPEQI5Z+0RjBUoS2
01xeeO+LJ6QPCi4p6ftYE6ZO4VJzUe2wzcKf9gpC6lXu1xh52D80MQNpBR+nNaq9
jEZzVImmFLI6lcYjCWuI26XGYadJF3mbUvhJVkDiVKz0CFK06bRgHyo1XOo9t/9M
Kk8EjyIvadPyHx2UlVk+W4UoIbP1k/4hkYvEhnEYIK067lwVNzIKdNDmJFeXBmo1
4jD8XmP2qoQQVKvfVk7FWY8tobcP8i/4vEwWe7zum42B/KGSic5lqXfQxwKlXY3a
LRo+KulHcduzK4xCUyooFM4AZVmQBwMkAJOwHX/LJ/t2ZxaUz76qXmjMxyFmvyAI
aD0Fj6CX1+uz3rbyH53LM9rf0tDuBeRBnk64EKAyrkBTr4rZKESmceq9lsuqYtNn
D5bFE2F7hM481b3tajYLI600lpkBrj5w5dnTZ+sFoK+zYndea07tibgoxoLNqzg3
FuGKtOz6TdXHvge0AyKXPMAniCkT87DLvKDBtUcCQiJuqVaUnAPfHLY41QImT9G7
tju+UOvnL2T8r5f5Vo6tiAj7/kWrMAj4KmqBmpWJG5Pstpkq6bynFRKSJsWomWqW
p+LTlIAbtDebd8dF25OpNQI6IvKCENvRKEy76Uaaq7lDxE6YB7HnXZCVYYefd5k/
IxyEzB2iTIdmLQFqkCFqV91YvRrsYlMyGiQxFqGAGlhS8ToPndDoiJ8y5J9tXfPM
/FT8ujU52emBEjdH2qnPrFql08vTv2DPmCvVn065cnFCQWsJr9xlJpn4jFFl9waW
LyG2K6hiwmki5YSg6M9v443W4qkD08BzKc2aYOCTmKSXdMwOrEymTPfkJZGnkgYl
fZGVPFCd0QXA5itHnJlB2Tez4EHipgRgGwf1N6LfQnLEw7oKCufNSm8b+7GdPNH/
JWIGoMVJnFaeAEchAb2ZLcDHOyYC/HUEBvXs03Vd6BSVW9i+ul4o/64ghBaGA+to
8Blb+aDmTMtgPEqn1Mz0LBgm3Pu04equVkgI3ikXwqQkBUq8Fojfdzye0CKkWWeq
H2Yqto4APqzBkDz/ca0/NPS62JZaLj+UZhtmlraNAvEs/nBLGsS5MYuLo+yNEZNa
Xhv6+yzKzCa7S9cJWJloD5Eh2MZQVka/zPVFjgKPm+JF5f3+hRs+6ThOr8AU9KaP
cWzp5YsZhkjzpVob8YcqXr4AmgpbiRWPYEtyN/xQB4D6RR8BQem5LTAT30PKJ+e+
xYTAH08OABwUpY1NVHn0LBvIAltbixtCVRfwIiD/36NfSPCwb1v0PYiKPLL4tcJT
2g8US9LSQxxp/8O4wehdjhqyWuMkDbPzTfs81k6yeQwijZm0QgwSUnKU18h+CPQy
dfa0elZJOb8UDRo0FSehldPDwv6AT0HfJL6ATKa0f7GWUWpr0ZSIbPscvkDikppu
JeG9rlMbUOpLWbBFDe8wS36kiMntAxz1bouggODsPV+s0z8fcsEticcrjYdBYrtH
47Tm3VDTa8KDUfrbtexrIrduzEM8zCXgFMMEmufz9wIXWygbbi6WfBxAueQWpHPP
bYzPBW9EL6zLQggy5+yoU1RJdoakkP+TrW3+fXcA31eZvqGlLCbYN/V8yHrsVljP
rV4VQ+xRiFLRMNzYZgnUfO/UCd1XtqPlVaHUCdEo1ajb6Ge64SWraFjDCTbAbtgh
cnEJylLmEBhCGDt+joykVWmzpjbtvjhes0o0DnbY09qQgtqxF5CZduw1s8r3jRpF
xWsu6tRDc/EYpVD4MBRC1Si7cG6ZvE5eZT6EpMUgQSFHT2gbJWi14/QCu4J3UMG6
5XVT+K/g85VnWFyXP6N1esPSBREKRCTD3vs49yA6uuhkCre+E32cX7ly3Y/Rv0j7
eFBUdP8DHGzuLEYeTVyO3ZxiJEAdVieF78gZlnvtPMBRPMF/ra0BTAi0sc0yiDVJ
aSAvRI+d6WhqtQ1QWl9EyzHfzG/ew5hM2FL71W8OItLXbfJBtUCKNGXuOAqv2wY5
NNcxg9rARXGuqXwZG9JeEznhf2gbRGpPBUrThEoHVBHsTnUaNnqaTbdXGvEPyhEy
rpT6HUV1G2NeJPU4kF9LEDhvpi/dwvOxoUMqaDug1ItgwAYYYJm7LqMSmQHSA32U
Sul935FtC4jCSteMcHJgIAGVoRlEPoQpGF7dECAD66yaKcH8f36Z0KnwvYCJaOeP
krr8vRXwquUT5QtLJCr0c6plwclzi22J4S7tWRLOenQg9s4mjht9rvI+rLRuyPc5
EjQ2wxo8tP3XHzSVHuwJ7F3Yew3nqRonhgpnRUeS7FH4qTRTJwEZ5d16o32KsihK
nTTCkFtixrH1T+et8h1dEMu8PXjcupp5f+LXFOvXrEyBkJOV1H9X9qsvv2KR2P9z
QnVKopSsFX2Xkt1nY2CTZxLThyeCWh50LJmrlgKKUFkrM1YW4NeveLq3GEe2XhP1
A92kqFsYQxT3Ge1iqbaH7F/gts43JshHpgjtUg9ZY8Dzx/Lt28gOGWeXTOT59LBn
+BdJNQTFWYzJM9XgEvGzXmesxgxDPugyNTzhrnzHJvIRn5gXDMhyF7rg4T1qhQXk
YC0BTy0eVRgN2CJZbC6/kfco8U0k9b/LmKfx1IxDd38Sjamup4OKp6oEn5UcJuhn
WcGNOvTmHNa0tKtcJ8temwSsi4v/74pKIhNqKCHC5+HmRMLZeRaF69+xmPKgRLhH
INhxIrZgFA2Jp99cZ2vYHfBr1SlOoUNTJ3XaZ5dnXk3oPWGpnt14jkDoKJnTcn9L
PXlM+Dpr6uP4PhNRKYBWl4yNB0+WvuvWKlUospx353U=
//pragma protect end_data_block
//pragma protect digest_block
R+YfoTcOog7QrEbYFAQujkTggpw=
//pragma protect end_digest_block
//pragma protect end_protected
